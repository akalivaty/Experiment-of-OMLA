//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1245, new_n1246, new_n1247, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(KEYINPUT65), .B(KEYINPUT0), .Z(new_n213));
  XNOR2_X1  g0013(.A(new_n212), .B(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(G20), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  INV_X1    g0018(.A(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(new_n214), .A2(KEYINPUT66), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n220), .B1(KEYINPUT66), .B2(new_n214), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT67), .Z(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n206), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(KEYINPUT68), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n227), .A2(new_n228), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n210), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT1), .Z(new_n235));
  NAND2_X1  g0035(.A1(new_n222), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT69), .Z(G361));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT70), .B(KEYINPUT2), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G226), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G68), .Z(new_n250));
  XNOR2_X1  g0050(.A(G58), .B(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  NAND3_X1  g0053(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(new_n215), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT74), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(new_n216), .A3(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G20), .A2(G33), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n256), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G1), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G13), .A3(G20), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(new_n202), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n255), .B1(new_n265), .B2(G20), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n268), .B2(new_n202), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT75), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n269), .B(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n264), .A2(new_n271), .A3(KEYINPUT9), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT9), .ZN(new_n273));
  XNOR2_X1  g0073(.A(new_n269), .B(KEYINPUT75), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(new_n263), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n272), .A2(new_n275), .ZN(new_n276));
  AND2_X1   g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  OAI21_X1  g0077(.A(KEYINPUT73), .B1(new_n277), .B2(new_n215), .ZN(new_n278));
  AND2_X1   g0078(.A1(G1), .A2(G13), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT73), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  OAI21_X1  g0085(.A(KEYINPUT71), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT3), .ZN(new_n287));
  INV_X1    g0087(.A(G33), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT71), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n289), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND4_X1  g0093(.A1(new_n286), .A2(new_n292), .A3(G222), .A4(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT72), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n286), .A2(new_n292), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n296), .A2(new_n293), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n297), .A2(G223), .B1(G77), .B2(new_n296), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n283), .B1(new_n295), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  OAI21_X1  g0100(.A(G274), .B1(new_n277), .B2(new_n215), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n265), .B1(G41), .B2(G45), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n279), .A2(new_n281), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n304), .A2(new_n302), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n303), .B1(G226), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NOR3_X1   g0107(.A1(new_n299), .A2(new_n300), .A3(new_n307), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n276), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(G200), .B1(new_n299), .B2(new_n307), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n309), .B(new_n310), .C1(KEYINPUT77), .C2(KEYINPUT10), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n299), .A2(new_n307), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G190), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n313), .A2(new_n310), .A3(new_n275), .A4(new_n272), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n313), .A2(KEYINPUT77), .A3(new_n275), .A4(new_n272), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT10), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G179), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n312), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n264), .A2(new_n271), .ZN(new_n320));
  INV_X1    g0120(.A(G169), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(new_n299), .B2(new_n307), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n319), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n311), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n259), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n266), .ZN(new_n326));
  INV_X1    g0126(.A(new_n268), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n259), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G58), .ZN(new_n331));
  INV_X1    g0131(.A(G68), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(G20), .B1(new_n333), .B2(new_n201), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n261), .A2(G159), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT16), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT81), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n289), .A2(new_n216), .A3(new_n291), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT7), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g0142(.A1(new_n289), .A2(KEYINPUT7), .A3(new_n216), .A4(new_n291), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n339), .B1(new_n344), .B2(G68), .ZN(new_n345));
  AOI211_X1 g0145(.A(KEYINPUT81), .B(new_n332), .C1(new_n342), .C2(new_n343), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n338), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT82), .ZN(new_n348));
  NOR2_X1   g0148(.A1(new_n284), .A2(new_n285), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT7), .B1(new_n349), .B2(new_n216), .ZN(new_n350));
  INV_X1    g0150(.A(new_n343), .ZN(new_n351));
  OAI21_X1  g0151(.A(G68), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT81), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n344), .A2(new_n339), .A3(G68), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT82), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n356), .A3(new_n338), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n348), .A2(new_n357), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n334), .A2(new_n335), .ZN(new_n359));
  NOR3_X1   g0159(.A1(new_n284), .A2(new_n285), .A3(KEYINPUT71), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n290), .B1(new_n289), .B2(new_n291), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n216), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n351), .B1(new_n362), .B2(new_n341), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n359), .B1(new_n363), .B2(new_n332), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n256), .B1(new_n364), .B2(new_n337), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n330), .B1(new_n358), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n303), .B1(G232), .B2(new_n305), .ZN(new_n367));
  OR2_X1    g0167(.A1(G223), .A2(G1698), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(G226), .B2(new_n293), .ZN(new_n369));
  OAI22_X1  g0169(.A1(new_n369), .A2(new_n349), .B1(new_n288), .B2(new_n224), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n277), .A2(KEYINPUT73), .A3(new_n215), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n280), .B1(new_n279), .B2(new_n281), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n367), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n375), .A2(new_n318), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(G169), .B2(new_n375), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT18), .B1(new_n366), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n356), .B1(new_n355), .B2(new_n338), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n359), .A2(KEYINPUT16), .ZN(new_n380));
  AOI211_X1 g0180(.A(KEYINPUT82), .B(new_n380), .C1(new_n353), .C2(new_n354), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n365), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(G200), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n375), .A2(new_n383), .ZN(new_n384));
  AND2_X1   g0184(.A1(KEYINPUT83), .A2(G190), .ZN(new_n385));
  NOR2_X1   g0185(.A1(KEYINPUT83), .A2(G190), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n384), .B1(new_n375), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n382), .A2(new_n329), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT17), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n377), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT18), .ZN(new_n393));
  AOI21_X1  g0193(.A(G20), .B1(new_n286), .B2(new_n292), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n343), .B1(new_n394), .B2(KEYINPUT7), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n336), .B1(new_n395), .B2(G68), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n255), .B1(new_n396), .B2(KEYINPUT16), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n397), .B1(new_n357), .B2(new_n348), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n392), .B(new_n393), .C1(new_n398), .C2(new_n330), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n366), .A2(KEYINPUT17), .A3(new_n388), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n378), .A2(new_n391), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n224), .A2(KEYINPUT15), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT15), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G87), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n216), .A2(G33), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n261), .ZN(new_n409));
  INV_X1    g0209(.A(G77), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n257), .A2(new_n409), .B1(new_n216), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n255), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n266), .A2(G77), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n413), .B1(new_n268), .B2(G77), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OR2_X1    g0215(.A1(new_n415), .A2(KEYINPUT76), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(KEYINPUT76), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n283), .B1(new_n296), .B2(new_n207), .ZN(new_n418));
  MUX2_X1   g0218(.A(G232), .B(G238), .S(G1698), .Z(new_n419));
  OAI21_X1  g0219(.A(new_n418), .B1(new_n296), .B2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n303), .B1(G244), .B2(new_n305), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n416), .B(new_n417), .C1(new_n383), .C2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n422), .A2(new_n300), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n423), .A2(G169), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n428), .A2(new_n415), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G179), .B2(new_n422), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  NOR3_X1   g0231(.A1(new_n324), .A2(new_n401), .A3(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT14), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT13), .ZN(new_n434));
  MUX2_X1   g0234(.A(G226), .B(G232), .S(G1698), .Z(new_n435));
  NAND3_X1  g0235(.A1(new_n435), .A2(new_n286), .A3(new_n292), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G97), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n373), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT78), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n440), .B1(new_n301), .B2(new_n302), .ZN(new_n441));
  INV_X1    g0241(.A(G274), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n442), .B1(new_n279), .B2(new_n281), .ZN(new_n443));
  INV_X1    g0243(.A(new_n302), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(KEYINPUT78), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n304), .A2(G238), .A3(new_n302), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n441), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n434), .B1(new_n439), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n283), .B1(new_n436), .B2(new_n437), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n441), .A2(new_n445), .A3(new_n446), .ZN(new_n450));
  NOR3_X1   g0250(.A1(new_n449), .A2(new_n450), .A3(KEYINPUT13), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n433), .B(G169), .C1(new_n448), .C2(new_n451), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n439), .A2(new_n447), .A3(new_n434), .ZN(new_n453));
  OAI21_X1  g0253(.A(KEYINPUT13), .B1(new_n449), .B2(new_n450), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n453), .A2(G179), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n453), .A2(new_n454), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n433), .B1(new_n457), .B2(G169), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT79), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g0259(.A1(new_n448), .A2(new_n451), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT14), .B1(new_n460), .B2(new_n321), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT79), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n461), .A2(new_n462), .A3(new_n455), .A4(new_n452), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n459), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT12), .ZN(new_n465));
  INV_X1    g0265(.A(new_n266), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(new_n332), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n266), .A2(KEYINPUT12), .A3(G68), .ZN(new_n468));
  OAI22_X1  g0268(.A1(new_n327), .A2(new_n332), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n261), .A2(G50), .B1(G20), .B2(new_n332), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(new_n410), .B2(new_n407), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n471), .A2(KEYINPUT11), .A3(new_n255), .ZN(new_n472));
  AOI21_X1  g0272(.A(KEYINPUT11), .B1(new_n471), .B2(new_n255), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n469), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n464), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n475), .B1(new_n460), .B2(G190), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n457), .A2(G200), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n476), .A2(KEYINPUT80), .A3(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT80), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n474), .B1(new_n459), .B2(new_n463), .ZN(new_n482));
  INV_X1    g0282(.A(new_n479), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n432), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(G41), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(KEYINPUT84), .A3(KEYINPUT5), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT5), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT84), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n490), .B1(new_n491), .B2(G41), .ZN(new_n492));
  INV_X1    g0292(.A(G45), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(G1), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n443), .A2(new_n489), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n492), .A2(new_n489), .A3(new_n494), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n304), .ZN(new_n497));
  INV_X1    g0297(.A(G270), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n296), .A2(G303), .ZN(new_n500));
  INV_X1    g0300(.A(G264), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G1698), .ZN(new_n502));
  OAI221_X1 g0302(.A(new_n502), .B1(G257), .B2(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n499), .B1(new_n504), .B2(new_n373), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G116), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n466), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n265), .A2(G33), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n256), .A2(new_n266), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n508), .B1(new_n510), .B2(new_n507), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G283), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n512), .B(new_n216), .C1(G33), .C2(new_n206), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n513), .B(new_n255), .C1(new_n216), .C2(G116), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT20), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n506), .A2(new_n519), .A3(G169), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT21), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n505), .A2(new_n387), .ZN(new_n523));
  OAI211_X1 g0323(.A(new_n523), .B(new_n518), .C1(new_n383), .C2(new_n505), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT88), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n283), .B1(new_n500), .B2(new_n503), .ZN(new_n526));
  OAI211_X1 g0326(.A(KEYINPUT21), .B(G169), .C1(new_n526), .C2(new_n499), .ZN(new_n527));
  INV_X1    g0327(.A(new_n499), .ZN(new_n528));
  INV_X1    g0328(.A(G303), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n286), .B2(new_n292), .ZN(new_n530));
  INV_X1    g0330(.A(new_n503), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n373), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n528), .A2(new_n532), .A3(G179), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n525), .B1(new_n534), .B2(new_n519), .ZN(new_n535));
  AOI211_X1 g0335(.A(KEYINPUT88), .B(new_n518), .C1(new_n527), .C2(new_n533), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n522), .B(new_n524), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n363), .A2(new_n207), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT6), .ZN(new_n539));
  NOR3_X1   g0339(.A1(new_n539), .A2(new_n206), .A3(G107), .ZN(new_n540));
  XNOR2_X1  g0340(.A(G97), .B(G107), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI22_X1  g0342(.A1(new_n542), .A2(new_n216), .B1(new_n410), .B2(new_n409), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n255), .B1(new_n538), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n286), .A2(new_n292), .A3(G250), .A4(G1698), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT4), .ZN(new_n546));
  INV_X1    g0346(.A(G244), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n546), .A2(new_n547), .A3(G1698), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n286), .A2(new_n292), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n293), .A2(G244), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n546), .B1(new_n349), .B2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n545), .A2(new_n549), .A3(new_n512), .A4(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n373), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n495), .B1(new_n497), .B2(new_n226), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G200), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n266), .A2(G97), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n256), .A2(new_n266), .A3(new_n509), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n558), .B1(new_n559), .B2(G97), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n554), .B1(new_n552), .B2(new_n373), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G190), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n544), .A2(new_n557), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n543), .B1(new_n395), .B2(G107), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n560), .B1(new_n564), .B2(new_n256), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n556), .A2(new_n321), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n561), .A2(new_n318), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n547), .A2(G1698), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(G238), .B2(G1698), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n570), .A2(new_n349), .B1(new_n288), .B2(new_n507), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n571), .A2(new_n373), .B1(new_n443), .B2(new_n494), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT86), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n304), .A2(G250), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT85), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(new_n493), .B2(G1), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n265), .A2(KEYINPUT85), .A3(G45), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n573), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n225), .B1(new_n279), .B2(new_n281), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n580), .A2(KEYINPUT86), .A3(new_n577), .A4(new_n576), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n572), .A2(G179), .A3(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n572), .A2(new_n582), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(new_n584), .B2(new_n321), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT19), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n216), .B1(new_n437), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(G87), .B2(new_n208), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n216), .B(G68), .C1(new_n284), .C2(new_n285), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n586), .B1(new_n407), .B2(new_n206), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(new_n255), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n559), .A2(new_n405), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n406), .A2(new_n466), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  OR2_X1    g0395(.A1(new_n595), .A2(KEYINPUT87), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(KEYINPUT87), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n585), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n383), .B1(new_n572), .B2(new_n582), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n599), .B1(G190), .B2(new_n584), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n559), .A2(G87), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n592), .A2(new_n601), .A3(new_n594), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n563), .A2(new_n568), .A3(new_n598), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n226), .A2(G1698), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(G250), .B2(G1698), .ZN(new_n607));
  INV_X1    g0407(.A(G294), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n607), .A2(new_n349), .B1(new_n288), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(new_n373), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n496), .A2(G264), .A3(new_n304), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n495), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(G169), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(KEYINPUT89), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT89), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n496), .A2(new_n615), .A3(G264), .A4(new_n304), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n614), .A2(new_n616), .B1(new_n373), .B2(new_n609), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n495), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n613), .B1(new_n618), .B2(new_n318), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT24), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n216), .B(G87), .C1(new_n284), .C2(new_n285), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(KEYINPUT22), .ZN(new_n622));
  OR3_X1    g0422(.A1(new_n224), .A2(KEYINPUT22), .A3(G20), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n622), .B1(new_n296), .B2(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n288), .A2(new_n507), .A3(G20), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT23), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n626), .B1(new_n216), .B2(G107), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n625), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n620), .B1(new_n624), .B2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n624), .A2(new_n620), .A3(new_n629), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n256), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n466), .A2(KEYINPUT25), .A3(new_n207), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT25), .B1(new_n466), .B2(new_n207), .ZN(new_n636));
  OAI22_X1  g0436(.A1(new_n635), .A2(new_n636), .B1(new_n510), .B2(new_n207), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n619), .B1(new_n633), .B2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n632), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n255), .B1(new_n639), .B2(new_n630), .ZN(new_n640));
  INV_X1    g0440(.A(new_n637), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n612), .A2(G190), .ZN(new_n642));
  AOI21_X1  g0442(.A(G200), .B1(new_n617), .B2(new_n495), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n638), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n537), .A2(new_n605), .A3(new_n645), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n487), .A2(new_n646), .ZN(G372));
  INV_X1    g0447(.A(new_n323), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n378), .A2(new_n399), .ZN(new_n649));
  INV_X1    g0449(.A(new_n430), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n482), .B1(new_n479), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n391), .A2(new_n400), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n649), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n311), .A2(new_n317), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n648), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n598), .A2(new_n604), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n656), .A2(new_n657), .A3(new_n568), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT91), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n568), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g0460(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT91), .A4(new_n567), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n602), .A2(KEYINPUT90), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT90), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n592), .A2(new_n601), .A3(new_n663), .A4(new_n594), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  AOI22_X1  g0465(.A1(new_n600), .A2(new_n665), .B1(new_n585), .B2(new_n595), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n660), .A2(new_n661), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n658), .B1(new_n657), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n585), .A2(new_n595), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n534), .A2(new_n519), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n638), .A2(new_n522), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n666), .A2(new_n644), .A3(new_n568), .A4(new_n563), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n669), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n655), .B1(new_n486), .B2(new_n675), .ZN(G369));
  NAND2_X1  g0476(.A1(new_n522), .A2(new_n670), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n265), .A2(new_n216), .A3(G13), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(G343), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n518), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n677), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n686), .B1(new_n537), .B2(new_n685), .ZN(new_n687));
  AND2_X1   g0487(.A1(new_n687), .A2(G330), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n684), .B1(new_n640), .B2(new_n641), .ZN(new_n689));
  OAI22_X1  g0489(.A1(new_n645), .A2(new_n689), .B1(new_n638), .B2(new_n684), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n638), .A2(new_n683), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n535), .A2(new_n536), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n683), .B1(new_n693), .B2(new_n522), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n694), .A2(new_n638), .A3(new_n644), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n691), .A2(new_n692), .A3(new_n695), .ZN(G399));
  INV_X1    g0496(.A(new_n211), .ZN(new_n697));
  OR3_X1    g0497(.A1(new_n697), .A2(KEYINPUT92), .A3(G41), .ZN(new_n698));
  OAI21_X1  g0498(.A(KEYINPUT92), .B1(new_n697), .B2(G41), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n224), .A2(new_n206), .A3(new_n207), .A4(new_n507), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n701), .A2(new_n265), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n703), .B1(new_n219), .B2(new_n701), .ZN(new_n704));
  XOR2_X1   g0504(.A(new_n704), .B(KEYINPUT28), .Z(new_n705));
  OAI21_X1  g0505(.A(new_n684), .B1(new_n668), .B2(new_n674), .ZN(new_n706));
  XOR2_X1   g0506(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n673), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n638), .B(new_n522), .C1(new_n535), .C2(new_n536), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n657), .B1(new_n656), .B2(new_n568), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n667), .B2(new_n657), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n711), .A2(new_n713), .A3(new_n669), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(KEYINPUT29), .A3(new_n684), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n646), .A2(new_n684), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT94), .ZN(new_n717));
  AND3_X1   g0517(.A1(new_n572), .A2(new_n717), .A3(new_n582), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n717), .B1(new_n572), .B2(new_n582), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n505), .A2(G179), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n720), .A2(new_n618), .A3(new_n556), .A4(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n561), .A2(new_n505), .A3(G179), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT93), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n584), .A2(new_n724), .A3(new_n617), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n614), .A2(new_n616), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(new_n610), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n572), .A2(new_n582), .ZN(new_n728));
  OAI21_X1  g0528(.A(KEYINPUT93), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n723), .B1(new_n725), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n722), .B1(new_n730), .B2(KEYINPUT30), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n556), .A2(new_n533), .ZN(new_n732));
  NOR3_X1   g0532(.A1(new_n727), .A2(new_n728), .A3(KEYINPUT93), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n724), .B1(new_n584), .B2(new_n617), .ZN(new_n734));
  OAI211_X1 g0534(.A(KEYINPUT30), .B(new_n732), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  OAI211_X1 g0536(.A(KEYINPUT31), .B(new_n683), .C1(new_n731), .C2(new_n736), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n683), .B1(new_n731), .B2(new_n736), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT31), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n716), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  AOI22_X1  g0541(.A1(new_n708), .A2(new_n715), .B1(G330), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n705), .B1(new_n742), .B2(G1), .ZN(G364));
  INV_X1    g0543(.A(G13), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n265), .B1(new_n745), .B2(G45), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  OR3_X1    g0547(.A1(new_n701), .A2(KEYINPUT96), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT96), .B1(new_n701), .B2(new_n747), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n215), .B1(G20), .B2(new_n321), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n216), .A2(new_n318), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n383), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(new_n387), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT98), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  NOR3_X1   g0558(.A1(new_n300), .A2(G179), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n216), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n758), .A2(G326), .B1(G294), .B2(new_n761), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n762), .A2(KEYINPUT99), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(KEYINPUT99), .ZN(new_n764));
  INV_X1    g0564(.A(new_n387), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n765), .A2(G200), .A3(new_n754), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(G322), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n216), .A2(G179), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n769), .A2(G190), .A3(G200), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n767), .A2(new_n768), .B1(new_n529), .B2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G190), .A2(G200), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G329), .ZN(new_n775));
  INV_X1    g0575(.A(G311), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n753), .A2(new_n772), .ZN(new_n777));
  OAI211_X1 g0577(.A(new_n775), .B(new_n296), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  NOR3_X1   g0578(.A1(new_n754), .A2(new_n383), .A3(G190), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  XOR2_X1   g0580(.A(KEYINPUT33), .B(G317), .Z(new_n781));
  NAND3_X1  g0581(.A1(new_n769), .A2(new_n300), .A3(G200), .ZN(new_n782));
  INV_X1    g0582(.A(G283), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n780), .A2(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n771), .A2(new_n778), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n763), .A2(new_n764), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n782), .A2(new_n207), .ZN(new_n787));
  INV_X1    g0587(.A(new_n296), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n410), .B2(new_n777), .ZN(new_n789));
  INV_X1    g0589(.A(new_n756), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n787), .B(new_n789), .C1(G50), .C2(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(new_n766), .A2(G58), .B1(G97), .B2(new_n761), .ZN(new_n792));
  INV_X1    g0592(.A(new_n770), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n779), .A2(G68), .B1(G87), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G159), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n773), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT97), .B(KEYINPUT32), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n791), .A2(new_n792), .A3(new_n794), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n752), .B1(new_n786), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n751), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n296), .A2(new_n697), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n805), .A2(G355), .B1(new_n507), .B2(new_n697), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n252), .A2(new_n493), .ZN(new_n807));
  INV_X1    g0607(.A(new_n349), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n697), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(G45), .B2(new_n218), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n806), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n800), .B1(new_n804), .B2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n803), .ZN(new_n813));
  OR2_X1    g0613(.A1(new_n687), .A2(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n750), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n687), .B(G330), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(new_n750), .B2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT100), .ZN(G396));
  OAI22_X1  g0618(.A1(new_n767), .A2(new_n608), .B1(new_n529), .B2(new_n756), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G107), .B2(new_n793), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n777), .A2(new_n507), .B1(new_n773), .B2(new_n776), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n788), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n782), .A2(new_n224), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G97), .B2(new_n761), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n820), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n780), .A2(KEYINPUT101), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT101), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n779), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n825), .B1(G283), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(new_n777), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n779), .A2(G150), .B1(G159), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  XOR2_X1   g0634(.A(KEYINPUT102), .B(G143), .Z(new_n835));
  OAI221_X1 g0635(.A(new_n833), .B1(new_n834), .B2(new_n756), .C1(new_n767), .C2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  INV_X1    g0639(.A(G132), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n808), .B1(new_n773), .B2(new_n840), .C1(new_n332), .C2(new_n782), .ZN(new_n841));
  OAI22_X1  g0641(.A1(new_n760), .A2(new_n331), .B1(new_n770), .B2(new_n202), .ZN(new_n842));
  NOR4_X1   g0642(.A1(new_n838), .A2(new_n839), .A3(new_n841), .A4(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n751), .B1(new_n831), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n751), .A2(new_n801), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n750), .B1(new_n410), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n650), .A2(new_n684), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n415), .A2(new_n684), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n426), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n847), .B1(new_n849), .B2(new_n650), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n844), .B(new_n846), .C1(new_n851), .C2(new_n802), .ZN(new_n852));
  INV_X1    g0652(.A(new_n750), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n706), .A2(new_n850), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n427), .A2(new_n430), .A3(new_n684), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n668), .B2(new_n674), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n741), .A2(G330), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n853), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n858), .A2(new_n859), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n852), .B1(new_n861), .B2(new_n862), .ZN(G384));
  NOR2_X1   g0663(.A1(new_n745), .A2(new_n265), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n336), .B1(new_n353), .B2(new_n354), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n255), .B1(new_n865), .B2(KEYINPUT16), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n866), .A2(KEYINPUT106), .B1(new_n357), .B2(new_n348), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT106), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n868), .B(new_n255), .C1(new_n865), .C2(KEYINPUT16), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n330), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n389), .B1(new_n870), .B2(new_n377), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n681), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT37), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n382), .A2(new_n329), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n392), .ZN(new_n875));
  INV_X1    g0675(.A(new_n681), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n875), .A2(new_n877), .A3(new_n878), .A4(new_n389), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n401), .A2(KEYINPUT107), .A3(new_n872), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT107), .B1(new_n401), .B2(new_n872), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n880), .B(KEYINPUT38), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n401), .A2(new_n872), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT107), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n401), .A2(KEYINPUT107), .A3(new_n872), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT38), .B1(new_n889), .B2(new_n880), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n884), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT105), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n476), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n482), .A2(KEYINPUT105), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n474), .A2(new_n684), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n483), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n893), .A2(new_n894), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n459), .A2(new_n463), .A3(new_n479), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n895), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n646), .A2(new_n684), .B1(new_n739), .B2(new_n738), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n850), .B1(new_n901), .B2(new_n737), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT40), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n482), .A2(KEYINPUT105), .ZN(new_n905));
  AOI211_X1 g0705(.A(new_n892), .B(new_n474), .C1(new_n459), .C2(new_n463), .ZN(new_n906));
  INV_X1    g0706(.A(new_n896), .ZN(new_n907));
  NOR3_X1   g0707(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n899), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n741), .B(new_n851), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT38), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n875), .A2(new_n877), .A3(new_n389), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n912), .B(new_n878), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n401), .A2(new_n874), .A3(new_n876), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n911), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n910), .B1(new_n883), .B2(new_n915), .ZN(new_n916));
  OAI22_X1  g0716(.A1(new_n891), .A2(new_n904), .B1(new_n916), .B2(new_n903), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n917), .A2(new_n487), .A3(new_n741), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(G330), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n917), .B1(new_n487), .B2(new_n741), .ZN(new_n920));
  OR2_X1    g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n883), .A2(new_n915), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(new_n911), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(KEYINPUT39), .A3(new_n883), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n893), .A2(new_n894), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(new_n684), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n924), .A2(new_n927), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n649), .A2(new_n876), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n926), .A2(new_n883), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n908), .A2(new_n909), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT104), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n857), .A2(new_n935), .A3(new_n847), .ZN(new_n936));
  INV_X1    g0736(.A(new_n669), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n709), .B2(new_n671), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n667), .A2(new_n657), .ZN(new_n939));
  OR3_X1    g0739(.A1(new_n656), .A2(new_n657), .A3(new_n568), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n855), .B1(new_n938), .B2(new_n941), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n430), .A2(new_n683), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT104), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n934), .B1(new_n936), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n932), .B1(new_n933), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n931), .A2(new_n946), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n708), .A2(new_n485), .A3(new_n432), .A4(new_n715), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n948), .A2(new_n655), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n947), .B(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n864), .B1(new_n921), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n950), .B2(new_n921), .ZN(new_n952));
  INV_X1    g0752(.A(new_n542), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n953), .A2(KEYINPUT35), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(KEYINPUT35), .ZN(new_n955));
  NAND4_X1  g0755(.A1(new_n954), .A2(G116), .A3(new_n217), .A4(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT36), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n333), .A2(new_n218), .A3(new_n410), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n958), .A2(KEYINPUT103), .B1(new_n202), .B2(G68), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(KEYINPUT103), .B2(new_n958), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(G1), .A3(new_n744), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n952), .A2(new_n957), .A3(new_n961), .ZN(G367));
  AND4_X1   g0762(.A1(new_n565), .A2(new_n566), .A3(new_n567), .A4(new_n683), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(KEYINPUT108), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n565), .A2(new_n683), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n563), .A2(new_n568), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n963), .A2(KEYINPUT108), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n691), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n970), .B(KEYINPUT109), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n665), .A2(new_n684), .ZN(new_n972));
  MUX2_X1   g0772(.A(new_n666), .B(new_n937), .S(new_n972), .Z(new_n973));
  NOR2_X1   g0773(.A1(new_n973), .A2(KEYINPUT43), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n971), .B(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n695), .A2(new_n969), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT42), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n568), .B1(new_n969), .B2(new_n638), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n977), .A2(KEYINPUT42), .B1(new_n684), .B2(new_n979), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n978), .A2(new_n980), .B1(KEYINPUT43), .B2(new_n973), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n975), .B(new_n981), .Z(new_n982));
  XNOR2_X1  g0782(.A(new_n700), .B(KEYINPUT41), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n695), .A2(new_n692), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n969), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT44), .Z(new_n986));
  NOR2_X1   g0786(.A1(new_n984), .A2(new_n969), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT45), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n986), .A2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(new_n691), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n695), .B1(new_n690), .B2(new_n694), .ZN(new_n991));
  XNOR2_X1  g0791(.A(new_n991), .B(new_n688), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n742), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n990), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n983), .B1(new_n995), .B2(new_n742), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n982), .B1(new_n996), .B2(new_n747), .ZN(new_n997));
  INV_X1    g0797(.A(new_n809), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n804), .B1(new_n211), .B2(new_n406), .C1(new_n245), .C2(new_n998), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n853), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n760), .A2(new_n332), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(G58), .B2(new_n793), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n782), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1003), .A2(G77), .ZN(new_n1004));
  INV_X1    g0804(.A(G150), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1002), .B(new_n1004), .C1(new_n767), .C2(new_n1005), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n777), .A2(new_n202), .B1(new_n773), .B2(new_n834), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n1006), .A2(new_n296), .A3(new_n1007), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n795), .B2(new_n829), .C1(new_n757), .C2(new_n835), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n1009), .B(KEYINPUT112), .Z(new_n1010));
  AND3_X1   g0810(.A1(new_n793), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n767), .A2(new_n529), .B1(new_n783), .B2(new_n777), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1011), .B(new_n1012), .C1(G107), .C2(new_n761), .ZN(new_n1013));
  AOI21_X1  g0813(.A(KEYINPUT46), .B1(new_n793), .B2(G116), .ZN(new_n1014));
  AOI22_X1  g0814(.A1(new_n830), .A2(G294), .B1(KEYINPUT110), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g0815(.A1(new_n1014), .A2(KEYINPUT110), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1016), .B1(new_n758), .B2(G311), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n808), .B1(new_n774), .B2(G317), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n206), .B2(new_n782), .ZN(new_n1019));
  XOR2_X1   g0819(.A(new_n1019), .B(KEYINPUT111), .Z(new_n1020));
  NAND4_X1  g0820(.A1(new_n1013), .A2(new_n1015), .A3(new_n1017), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1010), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT47), .Z(new_n1023));
  OAI221_X1 g0823(.A(new_n1000), .B1(new_n813), .B2(new_n973), .C1(new_n1023), .C2(new_n752), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n997), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT113), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(G387));
  AOI21_X1  g0827(.A(new_n808), .B1(new_n774), .B2(G326), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1028), .B1(new_n507), .B2(new_n782), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n829), .A2(new_n776), .B1(new_n757), .B2(new_n768), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT114), .ZN(new_n1031));
  OR2_X1    g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n766), .A2(G317), .B1(G303), .B2(new_n832), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT48), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n761), .A2(G283), .B1(new_n793), .B2(G294), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT49), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(KEYINPUT49), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1029), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n766), .A2(G50), .B1(G77), .B2(new_n793), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n795), .B2(new_n756), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n325), .A2(new_n780), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n808), .B1(new_n773), .B2(new_n1005), .C1(new_n332), .C2(new_n777), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n761), .A2(new_n405), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1048), .B1(new_n206), .B2(new_n782), .ZN(new_n1049));
  NOR4_X1   g0849(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .A4(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n751), .B1(new_n1043), .B2(new_n1050), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n242), .A2(new_n493), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n1052), .A2(new_n809), .B1(new_n702), .B2(new_n805), .ZN(new_n1053));
  AOI211_X1 g0853(.A(G45), .B(new_n702), .C1(G68), .C2(G77), .ZN(new_n1054));
  OR3_X1    g0854(.A1(new_n257), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1055));
  OAI21_X1  g0855(.A(KEYINPUT50), .B1(new_n257), .B2(G50), .ZN(new_n1056));
  AND3_X1   g0856(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n1053), .A2(new_n1057), .B1(G107), .B2(new_n211), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n750), .B1(new_n1058), .B2(new_n804), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1051), .B(new_n1059), .C1(new_n690), .C2(new_n813), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT115), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n994), .A2(new_n700), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n742), .B2(new_n992), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n992), .A2(new_n747), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1061), .A2(new_n1063), .A3(new_n1064), .ZN(G393));
  AOI21_X1  g0865(.A(new_n700), .B1(new_n990), .B2(new_n994), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(new_n994), .B2(new_n990), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n969), .A2(new_n803), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n1069), .A2(KEYINPUT116), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n1069), .A2(KEYINPUT116), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n804), .B1(new_n206), .B2(new_n211), .C1(new_n249), .C2(new_n998), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n853), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n830), .A2(G303), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(G294), .A2(new_n832), .B1(new_n774), .B2(G322), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n770), .A2(new_n783), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n787), .B(new_n1076), .C1(G116), .C2(new_n761), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1074), .A2(new_n296), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G317), .A2(new_n790), .B1(new_n766), .B2(G311), .ZN(new_n1079));
  XNOR2_X1  g0879(.A(new_n1079), .B(KEYINPUT52), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(G150), .A2(new_n790), .B1(new_n766), .B2(G159), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(new_n1081), .B(KEYINPUT51), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n808), .B1(new_n257), .B2(new_n777), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n835), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1083), .B1(new_n774), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n760), .A2(new_n410), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n823), .B(new_n1086), .C1(G68), .C2(new_n793), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1085), .B(new_n1087), .C1(new_n829), .C2(new_n202), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1078), .A2(new_n1080), .B1(new_n1082), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1073), .B1(new_n1089), .B2(new_n751), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1090), .B(KEYINPUT117), .ZN(new_n1091));
  NOR3_X1   g0891(.A1(new_n1070), .A2(new_n1071), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(new_n990), .B2(new_n747), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1067), .A2(new_n1093), .ZN(G390));
  NAND2_X1  g0894(.A1(new_n924), .A2(new_n927), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n944), .A2(new_n936), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n900), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n929), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n900), .A2(new_n902), .A3(G330), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n922), .A2(new_n929), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n714), .A2(new_n684), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n849), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n430), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n943), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n934), .ZN(new_n1106));
  OR2_X1    g0906(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1099), .A2(new_n1100), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1100), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n924), .A2(new_n927), .B1(new_n1097), .B2(new_n929), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1109), .B1(new_n1110), .B2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n432), .A2(new_n741), .A3(new_n485), .A4(G330), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n948), .A2(new_n655), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(KEYINPUT118), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT118), .ZN(new_n1116));
  NAND4_X1  g0916(.A1(new_n948), .A2(new_n655), .A3(new_n1116), .A4(new_n1113), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n741), .A2(new_n851), .A3(G330), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n934), .A2(new_n1119), .ZN(new_n1120));
  AND3_X1   g0920(.A1(new_n1120), .A2(new_n1100), .A3(new_n1105), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n1120), .A2(new_n1100), .B1(new_n936), .B2(new_n944), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1118), .A2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1108), .A2(new_n1112), .A3(new_n1124), .ZN(new_n1125));
  AND2_X1   g0925(.A1(new_n1125), .A2(new_n701), .ZN(new_n1126));
  INV_X1    g0926(.A(KEYINPUT119), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1127), .B(new_n1124), .C1(new_n1112), .C2(new_n1108), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1108), .A2(new_n1112), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1124), .ZN(new_n1130));
  AOI21_X1  g0930(.A(KEYINPUT119), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1126), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1108), .A2(new_n1112), .A3(new_n747), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1095), .A2(new_n801), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n750), .B1(new_n325), .B2(new_n845), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n782), .A2(new_n202), .ZN(new_n1136));
  OAI22_X1  g0936(.A1(new_n767), .A2(new_n840), .B1(new_n795), .B2(new_n760), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n1136), .B(new_n1137), .C1(G128), .C2(new_n790), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(KEYINPUT54), .B(G143), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n832), .A2(new_n1140), .B1(new_n774), .B2(G125), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT53), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1142), .B1(new_n770), .B2(new_n1005), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n793), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n830), .A2(G137), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1138), .A2(new_n788), .A3(new_n1141), .A4(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n767), .A2(new_n507), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1086), .B(new_n1147), .C1(G283), .C2(new_n790), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n830), .A2(G107), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n777), .A2(new_n206), .B1(new_n773), .B2(new_n608), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n788), .A2(new_n1150), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n793), .A2(G87), .B1(new_n1003), .B2(G68), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1148), .A2(new_n1149), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1146), .A2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1134), .B(new_n1135), .C1(new_n752), .C2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1132), .A2(new_n1133), .A3(new_n1155), .ZN(G378));
  INV_X1    g0956(.A(KEYINPUT122), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n947), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n931), .A2(new_n946), .A3(KEYINPUT122), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n320), .A2(new_n876), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n324), .B(new_n1160), .Z(new_n1161));
  XNOR2_X1  g0961(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1161), .B(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(new_n917), .B2(G330), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n910), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n903), .B1(new_n922), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n904), .B1(new_n926), .B2(new_n883), .ZN(new_n1168));
  OAI211_X1 g0968(.A(G330), .B(new_n1164), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n1158), .B(new_n1159), .C1(new_n1165), .C2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(G330), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1164), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1174), .A2(new_n931), .A3(new_n946), .A4(new_n1169), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1171), .A2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1118), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1125), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(KEYINPUT57), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(KEYINPUT123), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT123), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1171), .A2(new_n1175), .B1(new_n1125), .B2(new_n1177), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1182), .B2(KEYINPUT57), .ZN(new_n1183));
  INV_X1    g0983(.A(KEYINPUT57), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1184), .B1(new_n1125), .B2(new_n1177), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n947), .B1(new_n1165), .B2(new_n1170), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(new_n1175), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n700), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1180), .A2(new_n1183), .A3(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n750), .B1(new_n202), .B2(new_n845), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n808), .A2(G41), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1191), .B1(new_n783), .B2(new_n773), .C1(new_n406), .C2(new_n777), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1001), .B(new_n1192), .C1(G77), .C2(new_n793), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(new_n790), .A2(G116), .B1(G97), .B2(new_n779), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n766), .A2(G107), .B1(G58), .B2(new_n1003), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(new_n1196), .B(KEYINPUT120), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1197), .A2(KEYINPUT58), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1197), .A2(KEYINPUT58), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(G33), .A2(G41), .ZN(new_n1200));
  NOR3_X1   g1000(.A1(new_n1191), .A2(G50), .A3(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n790), .A2(G125), .B1(new_n793), .B2(new_n1140), .ZN(new_n1202));
  AOI22_X1  g1002(.A1(new_n766), .A2(G128), .B1(G132), .B2(new_n779), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n761), .A2(G150), .B1(new_n832), .B2(G137), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(KEYINPUT59), .ZN(new_n1207));
  INV_X1    g1007(.A(G124), .ZN(new_n1208));
  OAI221_X1 g1008(.A(new_n1200), .B1(new_n773), .B2(new_n1208), .C1(new_n795), .C2(new_n782), .ZN(new_n1209));
  XOR2_X1   g1009(.A(new_n1209), .B(KEYINPUT121), .Z(new_n1210));
  AND3_X1   g1010(.A1(new_n1206), .A2(new_n1207), .A3(new_n1210), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(new_n1198), .A2(new_n1199), .A3(new_n1201), .A4(new_n1211), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1190), .B1(new_n1212), .B2(new_n752), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1213), .B1(new_n1173), .B2(new_n801), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(new_n1176), .B2(new_n747), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1189), .A2(new_n1215), .ZN(G375));
  INV_X1    g1016(.A(new_n1123), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(new_n747), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G107), .A2(new_n832), .B1(new_n774), .B2(G303), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1219), .A2(new_n296), .A3(new_n1048), .A4(new_n1004), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n766), .A2(G283), .B1(G97), .B2(new_n793), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n608), .B2(new_n756), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1220), .B(new_n1222), .C1(G116), .C2(new_n830), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n829), .A2(new_n1139), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n761), .A2(G50), .B1(new_n793), .B2(G159), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n767), .B2(new_n834), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n349), .B1(new_n774), .B2(G128), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1005), .B2(new_n777), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n756), .A2(new_n840), .B1(new_n331), .B2(new_n782), .ZN(new_n1229));
  NOR4_X1   g1029(.A1(new_n1224), .A2(new_n1226), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n751), .B1(new_n1223), .B2(new_n1230), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n750), .B1(new_n332), .B2(new_n845), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1231), .B(new_n1232), .C1(new_n900), .C2(new_n802), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1218), .A2(new_n1233), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1177), .A2(new_n1217), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1124), .A2(new_n983), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1234), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(G381));
  INV_X1    g1039(.A(G375), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(G390), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1241));
  AND2_X1   g1041(.A1(new_n1241), .A2(new_n1238), .ZN(new_n1242));
  AND3_X1   g1042(.A1(new_n1132), .A2(new_n1133), .A3(new_n1155), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1240), .A2(new_n1026), .A3(new_n1242), .A4(new_n1243), .ZN(G407));
  NAND2_X1  g1044(.A1(new_n682), .A2(G213), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1247));
  OAI211_X1 g1047(.A(G407), .B(G213), .C1(G375), .C2(new_n1247), .ZN(G409));
  OAI21_X1  g1048(.A(new_n1188), .B1(new_n1179), .B2(KEYINPUT123), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1182), .A2(new_n1181), .A3(KEYINPUT57), .ZN(new_n1250));
  OAI211_X1 g1050(.A(G378), .B(new_n1215), .C1(new_n1249), .C2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n983), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1176), .A2(new_n1252), .A3(new_n1178), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1253), .A2(KEYINPUT124), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT124), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1182), .A2(new_n1255), .A3(new_n1252), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1214), .B1(new_n1187), .B2(new_n747), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1254), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1243), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1251), .A2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(new_n1245), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1124), .A2(new_n700), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1118), .A2(new_n1123), .A3(KEYINPUT60), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT125), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1266));
  OAI221_X1 g1066(.A(new_n1262), .B1(KEYINPUT60), .B2(new_n1235), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1234), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(G384), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1267), .A2(G384), .A3(new_n1268), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(G2897), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1245), .A2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1273), .A2(new_n1275), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1271), .B(new_n1272), .C1(new_n1274), .C2(new_n1245), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(KEYINPUT61), .B1(new_n1261), .B2(new_n1279), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1281), .B1(new_n1261), .B2(new_n1273), .ZN(new_n1282));
  INV_X1    g1082(.A(G390), .ZN(new_n1283));
  XOR2_X1   g1083(.A(G393), .B(G396), .Z(new_n1284));
  OAI21_X1  g1084(.A(new_n1283), .B1(new_n1284), .B2(KEYINPUT113), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1284), .A2(new_n1283), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1285), .A2(new_n1286), .A3(new_n1025), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1025), .B1(new_n1286), .B2(new_n1285), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1246), .B1(new_n1251), .B2(new_n1259), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1273), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1290), .A2(KEYINPUT63), .A3(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1280), .A2(new_n1282), .A3(new_n1289), .A4(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT62), .ZN(new_n1294));
  AND3_X1   g1094(.A1(new_n1290), .A2(new_n1294), .A3(new_n1291), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1296), .B1(new_n1290), .B2(new_n1278), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1294), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1298));
  NOR3_X1   g1098(.A1(new_n1295), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1293), .B1(new_n1299), .B2(new_n1289), .ZN(G405));
  OAI21_X1  g1100(.A(new_n1273), .B1(new_n1240), .B2(G378), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1251), .A2(KEYINPUT127), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(G375), .A2(new_n1291), .A3(new_n1243), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1301), .A2(new_n1302), .A3(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1302), .ZN(new_n1305));
  AND3_X1   g1105(.A1(G375), .A2(new_n1291), .A3(new_n1243), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1291), .B1(G375), .B2(new_n1243), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1305), .B1(new_n1306), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1304), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(new_n1289), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1304), .A2(new_n1308), .A3(new_n1289), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(G402));
endmodule


