//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 0 1 1 0 0 1 0 1 0 0 1 1 0 0 1 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:14 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n932,
    new_n933;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G57gat), .B(G85gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  NAND2_X1  g005(.A1(G155gat), .A2(G162gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT2), .ZN(new_n208));
  INV_X1    g007(.A(G141gat), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n209), .A2(G148gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n209), .A2(G148gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n208), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AND2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT78), .ZN(new_n215));
  NOR3_X1   g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G155gat), .ZN(new_n217));
  INV_X1    g016(.A(G162gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT78), .B1(new_n219), .B2(new_n207), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n212), .B1(new_n216), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT79), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n215), .B1(new_n213), .B2(new_n214), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n219), .A2(KEYINPUT78), .A3(new_n207), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT79), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n225), .A2(new_n226), .A3(new_n212), .ZN(new_n227));
  INV_X1    g026(.A(new_n210), .ZN(new_n228));
  XNOR2_X1  g027(.A(KEYINPUT80), .B(G148gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(new_n209), .ZN(new_n230));
  AOI22_X1  g029(.A1(KEYINPUT81), .A2(new_n208), .B1(new_n219), .B2(new_n207), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n208), .A2(KEYINPUT81), .ZN(new_n232));
  AND2_X1   g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI22_X1  g032(.A1(new_n222), .A2(new_n227), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(G127gat), .B(G134gat), .Z(new_n235));
  XNOR2_X1  g034(.A(G113gat), .B(G120gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n235), .B1(new_n236), .B2(KEYINPUT1), .ZN(new_n237));
  XOR2_X1   g036(.A(G113gat), .B(G120gat), .Z(new_n238));
  INV_X1    g037(.A(KEYINPUT1), .ZN(new_n239));
  XNOR2_X1  g038(.A(G127gat), .B(G134gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT4), .B1(new_n234), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT84), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n234), .A2(new_n244), .A3(new_n242), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n230), .A2(new_n232), .A3(new_n231), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n225), .A2(new_n226), .A3(new_n212), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n226), .B1(new_n225), .B2(new_n212), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n242), .B(new_n246), .C1(new_n247), .C2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT84), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n243), .B1(new_n251), .B2(KEYINPUT4), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n253), .B(new_n246), .C1(new_n247), .C2(new_n248), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT82), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n222), .A2(new_n227), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT82), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n256), .A2(new_n257), .A3(new_n253), .A4(new_n246), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n246), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n242), .B1(new_n260), .B2(KEYINPUT3), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n252), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G225gat), .A2(G233gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n206), .B1(new_n266), .B2(KEYINPUT39), .ZN(new_n267));
  OAI211_X1 g066(.A(new_n245), .B(new_n250), .C1(new_n234), .C2(new_n242), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT39), .B1(new_n268), .B2(new_n265), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n269), .B1(new_n263), .B2(new_n265), .ZN(new_n270));
  OAI21_X1  g069(.A(KEYINPUT90), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(KEYINPUT40), .ZN(new_n272));
  INV_X1    g071(.A(new_n206), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n274), .B1(new_n268), .B2(new_n265), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n265), .B1(new_n259), .B2(new_n261), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT4), .B1(new_n245), .B2(new_n250), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n249), .A2(KEYINPUT4), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT83), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n249), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n277), .B1(new_n278), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT85), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT85), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n277), .B(new_n286), .C1(new_n278), .C2(new_n283), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n276), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n252), .A2(new_n274), .A3(new_n277), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n273), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT40), .ZN(new_n292));
  OAI211_X1 g091(.A(KEYINPUT90), .B(new_n292), .C1(new_n267), .C2(new_n270), .ZN(new_n293));
  INV_X1    g092(.A(G183gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT27), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT27), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G183gat), .ZN(new_n297));
  INV_X1    g096(.A(G190gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT68), .ZN(new_n300));
  XOR2_X1   g099(.A(KEYINPUT69), .B(KEYINPUT28), .Z(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n301), .A2(new_n299), .A3(KEYINPUT68), .ZN(new_n304));
  INV_X1    g103(.A(G169gat), .ZN(new_n305));
  INV_X1    g104(.A(G176gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT26), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT26), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(G169gat), .B2(G176gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(G169gat), .A2(G176gat), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n310), .A2(new_n311), .B1(G183gat), .B2(G190gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n303), .A2(new_n304), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n315), .B(new_n316), .C1(G183gat), .C2(G190gat), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g119(.A(KEYINPUT66), .B(KEYINPUT23), .C1(G169gat), .C2(G176gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n311), .B(KEYINPUT67), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n317), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT25), .ZN(new_n325));
  OR3_X1    g124(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n314), .A2(KEYINPUT64), .ZN(new_n329));
  NOR2_X1   g128(.A1(new_n314), .A2(KEYINPUT64), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n328), .B(new_n316), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n311), .ZN(new_n332));
  AOI211_X1 g131(.A(KEYINPUT25), .B(new_n332), .C1(new_n320), .C2(new_n321), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n313), .A2(new_n325), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G226gat), .A2(G233gat), .ZN(new_n338));
  XOR2_X1   g137(.A(new_n338), .B(KEYINPUT75), .Z(new_n339));
  AOI22_X1  g138(.A1(new_n337), .A2(new_n338), .B1(new_n339), .B2(new_n335), .ZN(new_n340));
  XOR2_X1   g139(.A(G211gat), .B(G218gat), .Z(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT73), .ZN(new_n342));
  XNOR2_X1  g141(.A(G197gat), .B(G204gat), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT22), .ZN(new_n344));
  INV_X1    g143(.A(G211gat), .ZN(new_n345));
  INV_X1    g144(.A(G218gat), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n342), .B(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT74), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n340), .A2(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(new_n349), .B(KEYINPUT74), .Z(new_n352));
  AOI22_X1  g151(.A1(KEYINPUT25), .A2(new_n324), .B1(new_n331), .B2(new_n333), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n338), .B1(new_n353), .B2(new_n313), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n339), .B1(new_n335), .B2(new_n336), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n352), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT76), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT76), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n351), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G8gat), .B(G36gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G64gat), .B(G92gat), .ZN(new_n363));
  XOR2_X1   g162(.A(new_n362), .B(new_n363), .Z(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n356), .A3(new_n364), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT30), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(KEYINPUT77), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(KEYINPUT77), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT30), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n366), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n272), .A2(new_n291), .A3(new_n293), .A4(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(G78gat), .B(G106gat), .ZN(new_n374));
  INV_X1    g173(.A(G50gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n374), .B(new_n375), .ZN(new_n376));
  XNOR2_X1  g175(.A(KEYINPUT87), .B(KEYINPUT31), .ZN(new_n377));
  XNOR2_X1  g176(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n350), .B1(new_n259), .B2(new_n336), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT89), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(KEYINPUT29), .B1(new_n255), .B2(new_n258), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT89), .B1(new_n383), .B2(new_n350), .ZN(new_n384));
  INV_X1    g183(.A(G228gat), .ZN(new_n385));
  INV_X1    g184(.A(G233gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n253), .B1(new_n349), .B2(KEYINPUT29), .ZN(new_n387));
  AOI211_X1 g186(.A(new_n385), .B(new_n386), .C1(new_n387), .C2(new_n260), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n382), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G22gat), .ZN(new_n390));
  INV_X1    g189(.A(new_n348), .ZN(new_n391));
  OR2_X1    g190(.A1(new_n391), .A2(new_n341), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n341), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n392), .A2(new_n336), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT88), .ZN(new_n395));
  OR2_X1    g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT3), .B1(new_n394), .B2(new_n395), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n234), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI22_X1  g197(.A1(new_n380), .A2(new_n398), .B1(new_n385), .B2(new_n386), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n389), .A2(new_n390), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n390), .B1(new_n389), .B2(new_n399), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n379), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n389), .A2(new_n399), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(G22gat), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n389), .A2(new_n390), .A3(new_n399), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n378), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n373), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n287), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n249), .A2(KEYINPUT83), .A3(KEYINPUT4), .ZN(new_n411));
  AOI21_X1  g210(.A(KEYINPUT83), .B1(new_n249), .B2(KEYINPUT4), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT4), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n244), .B1(new_n234), .B2(new_n242), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n249), .A2(KEYINPUT84), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n286), .B1(new_n418), .B2(new_n277), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n275), .B1(new_n410), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n206), .A3(new_n289), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT6), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n291), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT91), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT94), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n355), .A2(new_n354), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n350), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT92), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT92), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n429), .A3(new_n350), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n428), .B(new_n430), .C1(new_n350), .C2(new_n340), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT37), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT38), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT93), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n435), .B1(new_n357), .B2(KEYINPUT37), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT37), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n351), .A2(new_n356), .A3(KEYINPUT93), .A4(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n436), .A2(new_n365), .A3(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n425), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(KEYINPUT38), .B1(new_n431), .B2(KEYINPUT37), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n438), .A2(new_n365), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n441), .A2(KEYINPUT94), .A3(new_n436), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(KEYINPUT6), .B(new_n273), .C1(new_n288), .C2(new_n290), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n437), .B1(new_n358), .B2(new_n360), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT38), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n445), .A2(new_n447), .A3(new_n367), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT91), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n291), .A2(new_n421), .A3(new_n449), .A4(new_n422), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n424), .A2(new_n444), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n409), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT70), .ZN(new_n453));
  INV_X1    g252(.A(new_n242), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n335), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n353), .A2(new_n242), .A3(new_n313), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(G227gat), .ZN(new_n458));
  NOR2_X1   g257(.A1(new_n458), .A2(new_n386), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n453), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n459), .ZN(new_n461));
  AOI211_X1 g260(.A(KEYINPUT70), .B(new_n461), .C1(new_n455), .C2(new_n456), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT32), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT33), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n464), .B1(new_n460), .B2(new_n462), .ZN(new_n465));
  XOR2_X1   g264(.A(G15gat), .B(G43gat), .Z(new_n466));
  XNOR2_X1  g265(.A(G71gat), .B(G99gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n463), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  OAI221_X1 g269(.A(KEYINPUT32), .B1(new_n464), .B2(new_n470), .C1(new_n460), .C2(new_n462), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n461), .ZN(new_n472));
  NAND2_X1  g271(.A1(KEYINPUT71), .A2(KEYINPUT34), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OR2_X1    g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(KEYINPUT71), .A2(KEYINPUT34), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n472), .B1(new_n476), .B2(new_n474), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n469), .A2(new_n471), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n469), .B2(new_n471), .ZN(new_n481));
  NOR3_X1   g280(.A1(new_n480), .A2(new_n481), .A3(KEYINPUT36), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n469), .A2(new_n471), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT72), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI211_X1 g284(.A(KEYINPUT72), .B(new_n478), .C1(new_n469), .C2(new_n471), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n482), .B1(new_n487), .B2(KEYINPUT36), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n423), .A2(new_n445), .ZN(new_n489));
  INV_X1    g288(.A(new_n372), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n488), .B1(new_n491), .B2(new_n407), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n489), .A2(new_n408), .A3(new_n490), .A4(new_n487), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(KEYINPUT35), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n424), .A2(new_n445), .A3(new_n450), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n480), .A2(new_n481), .ZN(new_n496));
  NOR4_X1   g295(.A1(new_n407), .A2(new_n496), .A3(KEYINPUT35), .A4(new_n372), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  AOI22_X1  g297(.A1(new_n452), .A2(new_n492), .B1(new_n494), .B2(new_n498), .ZN(new_n499));
  XNOR2_X1  g298(.A(G113gat), .B(G141gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(KEYINPUT95), .B(KEYINPUT11), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G169gat), .B(G197gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT12), .ZN(new_n505));
  XNOR2_X1  g304(.A(G15gat), .B(G22gat), .ZN(new_n506));
  INV_X1    g305(.A(G1gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT16), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(G1gat), .B2(new_n506), .ZN(new_n510));
  INV_X1    g309(.A(G8gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n375), .A2(G43gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(KEYINPUT97), .ZN(new_n515));
  XNOR2_X1  g314(.A(G43gat), .B(G50gat), .ZN(new_n516));
  OR2_X1    g315(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n518));
  AOI21_X1  g317(.A(G36gat), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G29gat), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n520), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n515), .B(new_n516), .C1(new_n519), .C2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n515), .B1(new_n519), .B2(new_n521), .ZN(new_n524));
  INV_X1    g323(.A(new_n516), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR3_X1    g325(.A1(new_n519), .A2(KEYINPUT15), .A3(new_n521), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n512), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT17), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n528), .B2(new_n523), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT17), .A4(new_n522), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n529), .B1(new_n533), .B2(new_n512), .ZN(new_n534));
  NAND2_X1  g333(.A1(G229gat), .A2(G233gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT98), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(KEYINPUT18), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  XOR2_X1   g338(.A(new_n535), .B(KEYINPUT13), .Z(new_n540));
  INV_X1    g339(.A(new_n512), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n528), .A2(new_n523), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n540), .B1(new_n543), .B2(new_n529), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n533), .A2(new_n512), .ZN(new_n545));
  INV_X1    g344(.A(new_n529), .ZN(new_n546));
  INV_X1    g345(.A(new_n538), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n535), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n539), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT96), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n505), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n548), .A2(new_n544), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n547), .B1(new_n534), .B2(new_n535), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n550), .B(new_n505), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n556), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n499), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT101), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(G155gat), .ZN(new_n561));
  XOR2_X1   g360(.A(G183gat), .B(G211gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT99), .B1(G71gat), .B2(G78gat), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NOR3_X1   g366(.A1(KEYINPUT99), .A2(G71gat), .A3(G78gat), .ZN(new_n568));
  OAI21_X1  g367(.A(new_n565), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT100), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(G57gat), .B(G64gat), .Z(new_n572));
  INV_X1    g371(.A(new_n565), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n572), .B1(KEYINPUT9), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(G71gat), .A2(G78gat), .ZN(new_n576));
  OR3_X1    g375(.A1(new_n574), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n578), .A2(KEYINPUT21), .ZN(new_n579));
  AND2_X1   g378(.A1(G231gat), .A2(G233gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n579), .B(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n581), .B(G127gat), .ZN(new_n582));
  INV_X1    g381(.A(new_n578), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT21), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n512), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n582), .A2(new_n585), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n564), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(new_n586), .A3(new_n563), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(KEYINPUT102), .A2(KEYINPUT7), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  NAND2_X1  g394(.A1(G99gat), .A2(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(G85gat), .ZN(new_n597));
  INV_X1    g396(.A(G92gat), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n596), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  AND2_X1   g398(.A1(new_n599), .A2(KEYINPUT103), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(KEYINPUT103), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n595), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(G99gat), .B(G106gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n603), .B(new_n595), .C1(new_n600), .C2(new_n601), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT104), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT105), .ZN(new_n609));
  OR2_X1    g408(.A1(new_n606), .A2(new_n607), .ZN(new_n610));
  AND3_X1   g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n609), .B1(new_n608), .B2(new_n610), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n542), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n610), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT105), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n533), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n613), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G190gat), .B(G218gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n613), .A2(new_n617), .A3(new_n622), .A4(new_n618), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(KEYINPUT106), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT107), .ZN(new_n626));
  XNOR2_X1  g425(.A(G134gat), .B(G162gat), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n625), .A2(new_n626), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n626), .B1(new_n625), .B2(new_n629), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n624), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n632), .ZN(new_n634));
  INV_X1    g433(.A(new_n624), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n634), .A2(new_n635), .A3(new_n630), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n592), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n583), .A2(new_n614), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n605), .A2(new_n606), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n578), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT10), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n578), .A2(KEYINPUT10), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n644), .B1(new_n615), .B2(new_n616), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n639), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n639), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n640), .A2(new_n642), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(G120gat), .B(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT108), .ZN(new_n651));
  XNOR2_X1  g450(.A(G176gat), .B(G204gat), .ZN(new_n652));
  XOR2_X1   g451(.A(new_n651), .B(new_n652), .Z(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n653), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n646), .A2(new_n648), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n558), .A2(new_n638), .A3(new_n658), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n659), .A2(new_n489), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n660), .B(new_n507), .ZN(G1324gat));
  INV_X1    g460(.A(KEYINPUT42), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n659), .A2(new_n490), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  AOI21_X1  g463(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(G8gat), .B1(new_n659), .B2(new_n490), .ZN(new_n666));
  INV_X1    g465(.A(new_n664), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n667), .B1(KEYINPUT109), .B2(new_n662), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n668), .B1(KEYINPUT109), .B2(new_n667), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n665), .A2(new_n666), .B1(new_n663), .B2(new_n669), .ZN(G1325gat));
  NAND2_X1  g469(.A1(new_n483), .A2(new_n484), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(new_n478), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n483), .A2(new_n484), .A3(new_n479), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(KEYINPUT36), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT36), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n496), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(G15gat), .B1(new_n659), .B2(new_n677), .ZN(new_n678));
  OR2_X1    g477(.A1(new_n496), .A2(G15gat), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n678), .B1(new_n659), .B2(new_n679), .ZN(G1326gat));
  NOR2_X1   g479(.A1(new_n659), .A2(new_n408), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  INV_X1    g482(.A(new_n637), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n499), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n589), .A2(new_n591), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n686), .A2(new_n557), .A3(new_n657), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT45), .ZN(new_n689));
  INV_X1    g488(.A(new_n489), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n520), .ZN(new_n691));
  OR3_X1    g490(.A1(new_n688), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(new_n499), .B2(new_n684), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n372), .B1(new_n423), .B2(new_n445), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n677), .B1(new_n695), .B2(new_n408), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n451), .B2(new_n409), .ZN(new_n697));
  AOI22_X1  g496(.A1(KEYINPUT35), .A2(new_n493), .B1(new_n495), .B2(new_n497), .ZN(new_n698));
  OAI211_X1 g497(.A(KEYINPUT44), .B(new_n637), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n694), .A2(new_n687), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n489), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n689), .B1(new_n688), .B2(new_n691), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n692), .A2(new_n701), .A3(new_n702), .ZN(G1328gat));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n704), .A2(KEYINPUT46), .ZN(new_n705));
  AOI21_X1  g504(.A(G36gat), .B1(new_n704), .B2(KEYINPUT46), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n372), .A2(new_n706), .ZN(new_n707));
  NOR4_X1   g506(.A1(new_n684), .A2(new_n686), .A3(new_n657), .A4(new_n707), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n558), .A2(new_n705), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n705), .B1(new_n558), .B2(new_n708), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(G36gat), .B1(new_n700), .B2(new_n490), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT111), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n711), .A2(new_n712), .A3(KEYINPUT111), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(G1329gat));
  OAI21_X1  g516(.A(G43gat), .B1(new_n700), .B2(new_n677), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n496), .A2(G43gat), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n685), .A2(new_n687), .A3(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT47), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n718), .A2(new_n720), .A3(KEYINPUT47), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(G1330gat));
  NAND4_X1  g524(.A1(new_n694), .A2(new_n407), .A3(new_n687), .A4(new_n699), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G50gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT112), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n685), .A2(new_n375), .A3(new_n407), .A4(new_n687), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n728), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n727), .B(new_n729), .C1(KEYINPUT112), .C2(KEYINPUT48), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(G1331gat));
  NAND2_X1  g533(.A1(new_n452), .A2(new_n492), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n494), .A2(new_n498), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT113), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n658), .A2(new_n556), .ZN(new_n739));
  NAND4_X1  g538(.A1(new_n737), .A2(new_n738), .A3(new_n638), .A4(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n638), .A2(new_n739), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT113), .B1(new_n499), .B2(new_n741), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n743), .A2(new_n690), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g544(.A1(new_n743), .A2(new_n372), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n747));
  XOR2_X1   g546(.A(KEYINPUT49), .B(G64gat), .Z(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n746), .B2(new_n748), .ZN(G1333gat));
  NAND3_X1  g548(.A1(new_n740), .A2(new_n742), .A3(new_n488), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(G71gat), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n496), .A2(G71gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n740), .A2(new_n742), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g552(.A(KEYINPUT114), .B(KEYINPUT50), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n751), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n754), .B1(new_n751), .B2(new_n753), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(G1334gat));
  NAND2_X1  g556(.A1(new_n743), .A2(new_n407), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT115), .B(G78gat), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1335gat));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n737), .A2(new_n637), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n686), .A2(new_n556), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n761), .B1(new_n762), .B2(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n685), .A2(KEYINPUT51), .A3(new_n763), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT116), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT116), .B(new_n761), .C1(new_n762), .C2(new_n764), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n489), .A2(G85gat), .A3(new_n658), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n764), .A2(new_n658), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n694), .A2(new_n699), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(G85gat), .B1(new_n773), .B2(new_n489), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n771), .A2(new_n774), .ZN(G1336gat));
  NOR3_X1   g574(.A1(new_n490), .A2(new_n658), .A3(G92gat), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n768), .A2(new_n769), .A3(new_n776), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n694), .A2(new_n372), .A3(new_n699), .A4(new_n772), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G92gat), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n776), .B(KEYINPUT117), .Z(new_n783));
  AOI22_X1  g582(.A1(new_n782), .A2(new_n783), .B1(new_n778), .B2(G92gat), .ZN(new_n784));
  OAI22_X1  g583(.A1(new_n777), .A2(new_n781), .B1(new_n784), .B2(new_n780), .ZN(G1337gat));
  NOR3_X1   g584(.A1(new_n496), .A2(new_n658), .A3(G99gat), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n768), .A2(new_n769), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(G99gat), .B1(new_n773), .B2(new_n677), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(G1338gat));
  NOR3_X1   g588(.A1(new_n408), .A2(G106gat), .A3(new_n658), .ZN(new_n790));
  AND3_X1   g589(.A1(new_n768), .A2(new_n769), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n694), .A2(new_n407), .A3(new_n699), .A4(new_n772), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G106gat), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n782), .A2(new_n790), .B1(new_n792), .B2(G106gat), .ZN(new_n796));
  OAI22_X1  g595(.A1(new_n791), .A2(new_n795), .B1(new_n796), .B2(new_n794), .ZN(G1339gat));
  INV_X1    g596(.A(KEYINPUT10), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n578), .B1(new_n610), .B2(new_n608), .ZN(new_n799));
  AND2_X1   g598(.A1(new_n578), .A2(new_n641), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI211_X1 g600(.A(KEYINPUT10), .B(new_n578), .C1(new_n611), .C2(new_n612), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n647), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n655), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n801), .A2(new_n802), .A3(new_n647), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n646), .A2(KEYINPUT54), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n805), .A2(new_n807), .A3(KEYINPUT55), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n556), .A2(new_n810), .A3(new_n656), .A4(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n813));
  OR3_X1    g612(.A1(new_n534), .A2(new_n813), .A3(new_n535), .ZN(new_n814));
  OR3_X1    g613(.A1(new_n543), .A2(new_n529), .A3(new_n540), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n534), .B2(new_n535), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n814), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n552), .A2(new_n553), .ZN(new_n818));
  AOI22_X1  g617(.A1(new_n817), .A2(new_n504), .B1(new_n818), .B2(new_n505), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n657), .A2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n812), .A2(new_n636), .A3(new_n633), .A4(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n810), .A2(new_n656), .A3(new_n811), .A4(new_n819), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n637), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n821), .A2(new_n592), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n684), .A2(new_n686), .A3(new_n557), .A4(new_n658), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n489), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n407), .A2(new_n485), .A3(new_n486), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n828), .A2(new_n490), .ZN(new_n829));
  AOI21_X1  g628(.A(G113gat), .B1(new_n829), .B2(new_n556), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n407), .B1(new_n824), .B2(new_n825), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n489), .A2(new_n372), .A3(new_n496), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n556), .A2(G113gat), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n830), .B1(new_n833), .B2(new_n834), .ZN(G1340gat));
  AOI21_X1  g634(.A(G120gat), .B1(new_n829), .B2(new_n657), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n657), .A2(G120gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n833), .B2(new_n837), .ZN(G1341gat));
  NAND3_X1  g637(.A1(new_n833), .A2(G127gat), .A3(new_n686), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n826), .A2(new_n490), .A3(new_n827), .A4(new_n686), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(G127gat), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n843), .B1(new_n840), .B2(new_n841), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n839), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT120), .ZN(G1342gat));
  AND2_X1   g645(.A1(new_n833), .A2(new_n637), .ZN(new_n847));
  INV_X1    g646(.A(G134gat), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n684), .A2(new_n372), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n828), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(KEYINPUT56), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n852), .B1(KEYINPUT56), .B2(new_n851), .ZN(G1343gat));
  NAND2_X1  g652(.A1(new_n824), .A2(new_n825), .ZN(new_n854));
  AND4_X1   g653(.A1(new_n690), .A2(new_n854), .A3(new_n407), .A4(new_n677), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n490), .A3(new_n556), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n209), .ZN(new_n857));
  AOI21_X1  g656(.A(KEYINPUT57), .B1(new_n854), .B2(new_n407), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n859));
  AOI211_X1 g658(.A(new_n859), .B(new_n408), .C1(new_n824), .C2(new_n825), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NOR3_X1   g660(.A1(new_n488), .A2(new_n489), .A3(new_n372), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n556), .A2(G141gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n857), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT58), .ZN(new_n866));
  XNOR2_X1  g665(.A(new_n865), .B(new_n866), .ZN(G1344gat));
  INV_X1    g666(.A(new_n229), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n855), .A2(new_n868), .A3(new_n490), .A4(new_n657), .ZN(new_n869));
  XOR2_X1   g668(.A(new_n869), .B(KEYINPUT121), .Z(new_n870));
  OAI211_X1 g669(.A(new_n657), .B(new_n862), .C1(new_n858), .C2(new_n860), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G148gat), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT59), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n868), .A2(KEYINPUT59), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT122), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n871), .A2(KEYINPUT122), .A3(new_n875), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n874), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n873), .B1(new_n872), .B2(KEYINPUT59), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n870), .B1(new_n880), .B2(new_n881), .ZN(G1345gat));
  OAI21_X1  g681(.A(G155gat), .B1(new_n863), .B2(new_n592), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n855), .A2(new_n217), .A3(new_n490), .A4(new_n686), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1346gat));
  NAND3_X1  g684(.A1(new_n855), .A2(new_n218), .A3(new_n850), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT124), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n863), .B2(new_n684), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(G162gat), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n863), .A2(new_n887), .A3(new_n684), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(G1347gat));
  NOR3_X1   g690(.A1(new_n690), .A2(new_n490), .A3(new_n496), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n831), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(new_n305), .A3(new_n557), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n690), .B1(new_n824), .B2(new_n825), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n895), .A2(new_n372), .A3(new_n827), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(new_n556), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n894), .B1(new_n897), .B2(new_n305), .ZN(G1348gat));
  NOR3_X1   g697(.A1(new_n893), .A2(new_n306), .A3(new_n658), .ZN(new_n899));
  AOI21_X1  g698(.A(G176gat), .B1(new_n896), .B2(new_n657), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n900), .A2(KEYINPUT125), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(KEYINPUT125), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(G1349gat));
  NAND4_X1  g702(.A1(new_n896), .A2(new_n295), .A3(new_n297), .A4(new_n686), .ZN(new_n904));
  OAI21_X1  g703(.A(G183gat), .B1(new_n893), .B2(new_n592), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n907));
  XOR2_X1   g706(.A(new_n906), .B(new_n907), .Z(G1350gat));
  NAND3_X1  g707(.A1(new_n896), .A2(new_n298), .A3(new_n637), .ZN(new_n909));
  OAI21_X1  g708(.A(G190gat), .B1(new_n893), .B2(new_n684), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n910), .A2(KEYINPUT61), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(KEYINPUT61), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n909), .B1(new_n911), .B2(new_n912), .ZN(G1351gat));
  XNOR2_X1  g712(.A(KEYINPUT127), .B(G197gat), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n488), .A2(new_n690), .A3(new_n490), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n861), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n914), .B1(new_n916), .B2(new_n557), .ZN(new_n917));
  AND4_X1   g716(.A1(new_n407), .A2(new_n895), .A3(new_n372), .A4(new_n677), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n557), .A2(new_n914), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n917), .A2(new_n920), .ZN(G1352gat));
  INV_X1    g720(.A(G204gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n918), .A2(new_n922), .A3(new_n657), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT62), .Z(new_n924));
  OAI21_X1  g723(.A(G204gat), .B1(new_n916), .B2(new_n658), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1353gat));
  NAND3_X1  g725(.A1(new_n918), .A2(new_n345), .A3(new_n686), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n861), .A2(new_n686), .A3(new_n915), .ZN(new_n928));
  AND3_X1   g727(.A1(new_n928), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT63), .B1(new_n928), .B2(G211gat), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n927), .B1(new_n929), .B2(new_n930), .ZN(G1354gat));
  OAI21_X1  g730(.A(G218gat), .B1(new_n916), .B2(new_n684), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n918), .A2(new_n346), .A3(new_n637), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(G1355gat));
endmodule


