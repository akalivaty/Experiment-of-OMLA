//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n551, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n618, new_n619, new_n622, new_n623, new_n625, new_n626,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1188;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XOR2_X1   g014(.A(KEYINPUT64), .B(G57), .Z(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XOR2_X1   g020(.A(new_n445), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT67), .ZN(new_n464));
  AND2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  AOI22_X1  g043(.A1(G101), .A2(new_n464), .B1(new_n468), .B2(G137), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  XNOR2_X1  g045(.A(new_n470), .B(KEYINPUT66), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OR2_X1    g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NAND2_X1  g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g050(.A(G2105), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n469), .A2(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n468), .A2(G136), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT68), .Z(new_n479));
  AOI21_X1  g054(.A(new_n462), .B1(new_n473), .B2(new_n474), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT69), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n479), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI211_X1 g061(.A(G138), .B(new_n462), .C1(new_n465), .C2(new_n466), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(new_n462), .A3(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT70), .B1(new_n467), .B2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n473), .A2(new_n474), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n493));
  AND3_X1   g068(.A1(new_n489), .A2(new_n462), .A3(G138), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n488), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G2105), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(G126), .B2(new_n480), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G62), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT72), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n505), .A2(new_n506), .B1(G75), .B2(G543), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n504), .A2(KEYINPUT72), .A3(G62), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n503), .B2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT6), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G651), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(G543), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n515), .A2(new_n504), .A3(new_n516), .ZN(new_n518));
  INV_X1    g093(.A(G88), .ZN(new_n519));
  OAI22_X1  g094(.A1(new_n510), .A2(new_n517), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n509), .A2(new_n520), .ZN(G166));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n524));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n523), .A2(new_n524), .B1(new_n504), .B2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  INV_X1    g102(.A(G51), .ZN(new_n528));
  OAI221_X1 g103(.A(new_n526), .B1(new_n518), .B2(new_n527), .C1(new_n528), .C2(new_n517), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AOI22_X1  g105(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n531), .A2(new_n503), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n517), .ZN(new_n535));
  INV_X1    g110(.A(new_n518), .ZN(new_n536));
  AOI22_X1  g111(.A1(G52), .A2(new_n535), .B1(new_n536), .B2(G90), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n534), .A2(new_n538), .ZN(G171));
  AOI22_X1  g114(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n503), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G43), .ZN(new_n543));
  INV_X1    g118(.A(G81), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n543), .A2(new_n517), .B1(new_n518), .B2(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n545), .A2(KEYINPUT74), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n542), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  AOI22_X1  g130(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n503), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(G78), .A2(G543), .ZN(new_n559));
  AND2_X1   g134(.A1(KEYINPUT5), .A2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(KEYINPUT5), .A2(G543), .ZN(new_n561));
  NOR2_X1   g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT75), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n558), .A2(new_n565), .B1(new_n536), .B2(G91), .ZN(new_n566));
  INV_X1    g141(.A(G53), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT9), .B1(new_n517), .B2(new_n567), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n511), .A2(new_n514), .B1(KEYINPUT6), .B2(new_n503), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n569), .A2(new_n570), .A3(G53), .A4(G543), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n566), .A2(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  OR2_X1    g149(.A1(new_n509), .A2(new_n520), .ZN(G303));
  NAND3_X1  g150(.A1(new_n569), .A2(G87), .A3(new_n504), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n569), .A2(G49), .A3(G543), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  OAI21_X1  g154(.A(G61), .B1(new_n560), .B2(new_n561), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g157(.A(KEYINPUT76), .B1(new_n582), .B2(G651), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  AOI211_X1 g159(.A(new_n584), .B(new_n503), .C1(new_n580), .C2(new_n581), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n569), .A2(G48), .A3(G543), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n569), .A2(G86), .A3(new_n504), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G305));
  AOI22_X1  g166(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  NOR2_X1   g167(.A1(new_n592), .A2(new_n503), .ZN(new_n593));
  XOR2_X1   g168(.A(new_n593), .B(KEYINPUT77), .Z(new_n594));
  NAND2_X1  g169(.A1(new_n536), .A2(G85), .ZN(new_n595));
  XOR2_X1   g170(.A(KEYINPUT78), .B(G47), .Z(new_n596));
  NAND2_X1  g171(.A1(new_n535), .A2(new_n596), .ZN(new_n597));
  AND3_X1   g172(.A1(new_n595), .A2(new_n597), .A3(KEYINPUT79), .ZN(new_n598));
  AOI21_X1  g173(.A(KEYINPUT79), .B1(new_n595), .B2(new_n597), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n594), .B1(new_n598), .B2(new_n599), .ZN(G290));
  INV_X1    g175(.A(G92), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n518), .A2(new_n601), .ZN(new_n602));
  OR2_X1    g177(.A1(new_n602), .A2(KEYINPUT10), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(KEYINPUT10), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(G79), .A2(G543), .ZN(new_n606));
  INV_X1    g181(.A(G66), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n562), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G651), .ZN(new_n609));
  INV_X1    g184(.A(G54), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n517), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n605), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n614), .B2(G171), .ZN(G284));
  OAI21_X1  g191(.A(new_n615), .B1(new_n614), .B2(G171), .ZN(G321));
  NAND2_X1  g192(.A1(G286), .A2(G868), .ZN(new_n618));
  INV_X1    g193(.A(G299), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G297));
  OAI21_X1  g195(.A(new_n618), .B1(new_n619), .B2(G868), .ZN(G280));
  AOI21_X1  g196(.A(new_n611), .B1(new_n603), .B2(new_n604), .ZN(new_n622));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n548), .A2(new_n614), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n613), .A2(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(new_n614), .ZN(G323));
  XNOR2_X1  g202(.A(KEYINPUT80), .B(KEYINPUT11), .ZN(new_n628));
  XNOR2_X1  g203(.A(G323), .B(new_n628), .ZN(G282));
  NAND2_X1  g204(.A1(new_n464), .A2(new_n492), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT12), .Z(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2100), .Z(new_n632));
  XOR2_X1   g207(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n468), .A2(G135), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n480), .A2(G123), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n462), .A2(G111), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  OAI211_X1 g214(.A(new_n636), .B(new_n637), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND3_X1  g216(.A1(new_n634), .A2(new_n635), .A3(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT82), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2427), .B(G2430), .Z(new_n646));
  OR2_X1    g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n646), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(KEYINPUT14), .A3(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G2451), .B(G2454), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1341), .B(G1348), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n649), .B(new_n653), .Z(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n654), .A2(new_n655), .ZN(new_n657));
  AND3_X1   g232(.A1(new_n656), .A2(G14), .A3(new_n657), .ZN(G401));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  XNOR2_X1  g234(.A(G2067), .B(G2678), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n661), .A2(KEYINPUT17), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n659), .A2(new_n660), .ZN(new_n663));
  AOI21_X1  g238(.A(KEYINPUT18), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2072), .B(G2078), .Z(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XNOR2_X1  g244(.A(G1971), .B(G1976), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1956), .B(G2474), .ZN(new_n673));
  XNOR2_X1  g248(.A(G1961), .B(G1966), .ZN(new_n674));
  NOR3_X1   g249(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n675), .B(KEYINPUT20), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n673), .A2(new_n674), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n672), .A2(KEYINPUT84), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n681), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n682), .A3(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT85), .Z(new_n685));
  XNOR2_X1  g260(.A(G1991), .B(G1996), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n685), .B(new_n690), .ZN(G229));
  NAND2_X1  g266(.A1(new_n468), .A2(G139), .ZN(new_n692));
  XOR2_X1   g267(.A(new_n692), .B(KEYINPUT90), .Z(new_n693));
  NAND3_X1  g268(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT25), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  AOI22_X1  g271(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n693), .B(new_n696), .C1(new_n462), .C2(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G33), .B(new_n698), .S(G29), .Z(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G2072), .ZN(new_n700));
  XOR2_X1   g275(.A(new_n700), .B(KEYINPUT91), .Z(new_n701));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G4), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(new_n622), .B2(new_n702), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n701), .B1(G1348), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT86), .B(G16), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n707), .A2(G19), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n549), .B2(new_n707), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(G1341), .Z(new_n710));
  OAI211_X1 g285(.A(new_n705), .B(new_n710), .C1(G1348), .C2(new_n704), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n699), .A2(G2072), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G27), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G164), .B2(new_n713), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(G2078), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT31), .B(G11), .Z(new_n718));
  XNOR2_X1  g293(.A(KEYINPUT30), .B(G28), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n718), .B1(new_n713), .B2(new_n719), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(new_n640), .B2(new_n713), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n713), .A2(G26), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n468), .A2(G140), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n480), .A2(G128), .ZN(new_n725));
  OR2_X1    g300(.A1(G104), .A2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n726), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n723), .B1(new_n729), .B2(new_n713), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n721), .B1(new_n730), .B2(G2067), .ZN(new_n731));
  INV_X1    g306(.A(G2084), .ZN(new_n732));
  NAND2_X1  g307(.A1(G160), .A2(G29), .ZN(new_n733));
  INV_X1    g308(.A(G34), .ZN(new_n734));
  AOI21_X1  g309(.A(G29), .B1(new_n734), .B2(KEYINPUT24), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(KEYINPUT24), .B2(new_n734), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n733), .A2(new_n736), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n731), .B1(G2067), .B2(new_n730), .C1(new_n732), .C2(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G171), .A2(new_n702), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G5), .B2(new_n702), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n738), .B1(new_n741), .B2(G1961), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n713), .A2(G32), .ZN(new_n743));
  AOI22_X1  g318(.A1(G105), .A2(new_n464), .B1(new_n468), .B2(G141), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n480), .A2(G129), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT26), .Z(new_n747));
  NAND3_X1  g322(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT92), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n748), .A2(new_n749), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n743), .B1(new_n753), .B2(new_n713), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT93), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n717), .B(new_n742), .C1(new_n755), .C2(new_n757), .ZN(new_n758));
  OAI21_X1  g333(.A(KEYINPUT94), .B1(G16), .B2(G21), .ZN(new_n759));
  NOR2_X1   g334(.A1(G286), .A2(new_n702), .ZN(new_n760));
  MUX2_X1   g335(.A(new_n759), .B(KEYINPUT94), .S(new_n760), .Z(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1966), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n713), .A2(G35), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n763), .B1(G162), .B2(new_n713), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT29), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n762), .B1(new_n765), .B2(G2090), .ZN(new_n766));
  NOR3_X1   g341(.A1(new_n711), .A2(new_n758), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n702), .A2(G23), .ZN(new_n768));
  INV_X1    g343(.A(G288), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n768), .B1(new_n769), .B2(new_n702), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT33), .ZN(new_n771));
  INV_X1    g346(.A(G1976), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n702), .A2(G6), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(new_n590), .B2(new_n702), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT32), .B(G1981), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT88), .ZN(new_n777));
  XOR2_X1   g352(.A(new_n775), .B(new_n777), .Z(new_n778));
  NOR2_X1   g353(.A1(new_n707), .A2(G22), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G166), .B2(new_n707), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT89), .B(G1971), .Z(new_n781));
  XOR2_X1   g356(.A(new_n780), .B(new_n781), .Z(new_n782));
  NOR3_X1   g357(.A1(new_n773), .A2(new_n778), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT87), .B(KEYINPUT34), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n468), .A2(G131), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n480), .A2(G119), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n462), .A2(G107), .ZN(new_n789));
  OAI21_X1  g364(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n787), .B(new_n788), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G25), .B(new_n791), .S(G29), .Z(new_n792));
  XOR2_X1   g367(.A(KEYINPUT35), .B(G1991), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  AND2_X1   g369(.A1(new_n706), .A2(G24), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G290), .B2(new_n707), .ZN(new_n796));
  INV_X1    g371(.A(G1986), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n797), .B2(new_n796), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n785), .A2(new_n786), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT36), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n755), .A2(new_n757), .ZN(new_n802));
  INV_X1    g377(.A(G1961), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n740), .A2(new_n803), .B1(new_n732), .B2(new_n737), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT95), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n765), .A2(G2090), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n706), .A2(G20), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT23), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n619), .B2(new_n702), .ZN(new_n812));
  INV_X1    g387(.A(G1956), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n809), .A2(new_n814), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n807), .B1(new_n808), .B2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n815), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n817), .A2(KEYINPUT96), .B1(new_n805), .B2(new_n806), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n767), .A2(new_n801), .A3(new_n816), .A4(new_n818), .ZN(G150));
  INV_X1    g394(.A(G150), .ZN(G311));
  NAND2_X1  g395(.A1(new_n535), .A2(G55), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n536), .A2(G93), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n823), .A2(new_n503), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(G860), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  NAND2_X1  g402(.A1(new_n622), .A2(G559), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(KEYINPUT97), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT38), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n548), .A2(new_n825), .ZN(new_n831));
  INV_X1    g406(.A(new_n825), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n832), .B(new_n542), .C1(new_n546), .C2(new_n547), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n830), .B(new_n834), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n835), .A2(KEYINPUT39), .ZN(new_n836));
  INV_X1    g411(.A(G860), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n835), .B2(KEYINPUT39), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n827), .B1(new_n836), .B2(new_n838), .ZN(G145));
  XNOR2_X1  g414(.A(new_n752), .B(new_n728), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n468), .A2(G142), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT98), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n843));
  INV_X1    g418(.A(G118), .ZN(new_n844));
  AOI22_X1  g419(.A1(new_n843), .A2(KEYINPUT99), .B1(new_n844), .B2(G2105), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(KEYINPUT99), .B2(new_n843), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n480), .A2(G130), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n842), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n840), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n698), .B(new_n501), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n631), .B(new_n791), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n849), .B(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(G160), .B(new_n640), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G162), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(G37), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n853), .A2(new_n855), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(G395));
  XNOR2_X1  g436(.A(new_n834), .B(new_n626), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT101), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n613), .A2(new_n863), .A3(new_n619), .ZN(new_n864));
  OAI21_X1  g439(.A(KEYINPUT101), .B1(new_n622), .B2(G299), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n622), .A2(G299), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  OR2_X1    g443(.A1(new_n862), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT41), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n867), .B(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n862), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT42), .ZN(new_n874));
  NAND2_X1  g449(.A1(G290), .A2(new_n769), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n594), .B(G288), .C1(new_n599), .C2(new_n598), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  NAND2_X1  g453(.A1(G303), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(G166), .A2(KEYINPUT102), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n879), .A2(G305), .A3(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(G305), .B1(new_n879), .B2(new_n880), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n877), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n885), .A2(new_n875), .A3(new_n876), .A4(new_n881), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n873), .A2(KEYINPUT42), .ZN(new_n889));
  AND3_X1   g464(.A1(new_n874), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n888), .B1(new_n874), .B2(new_n889), .ZN(new_n891));
  OAI21_X1  g466(.A(G868), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n892), .B1(G868), .B2(new_n832), .ZN(G295));
  OAI21_X1  g468(.A(new_n892), .B1(G868), .B2(new_n832), .ZN(G331));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT104), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n896), .B(G286), .C1(new_n534), .C2(new_n538), .ZN(new_n897));
  NAND2_X1  g472(.A1(G286), .A2(new_n896), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n532), .B(KEYINPUT73), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n536), .A2(G89), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n535), .A2(G51), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT104), .A4(new_n526), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n898), .A2(new_n899), .A3(new_n902), .A4(new_n537), .ZN(new_n903));
  AND2_X1   g478(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n904), .A2(KEYINPUT105), .A3(new_n831), .A4(new_n833), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n831), .A2(new_n833), .A3(new_n897), .A4(new_n903), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n897), .A2(new_n903), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n834), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n908), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n895), .B1(new_n911), .B2(new_n868), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n906), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n871), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g490(.A1(new_n911), .A2(new_n895), .A3(new_n868), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n887), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n913), .ZN(new_n918));
  AOI22_X1  g493(.A1(new_n871), .A2(new_n911), .B1(new_n918), .B2(new_n867), .ZN(new_n919));
  AOI21_X1  g494(.A(G37), .B1(new_n919), .B2(new_n888), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n917), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n871), .A2(new_n911), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(new_n867), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n888), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n857), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n919), .A2(new_n888), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT43), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n922), .A2(new_n928), .ZN(new_n929));
  XOR2_X1   g504(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(KEYINPUT107), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT107), .ZN(new_n933));
  AOI211_X1 g508(.A(new_n933), .B(new_n930), .C1(new_n922), .C2(new_n928), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n921), .B1(new_n917), .B2(new_n920), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n920), .B1(new_n888), .B2(new_n919), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT44), .B1(new_n936), .B2(KEYINPUT43), .ZN(new_n937));
  OAI22_X1  g512(.A1(new_n932), .A2(new_n934), .B1(new_n935), .B2(new_n937), .ZN(G397));
  INV_X1    g513(.A(G1384), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT45), .B1(new_n501), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n464), .A2(G101), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n468), .A2(G137), .ZN(new_n942));
  AND4_X1   g517(.A1(G40), .A2(new_n941), .A3(new_n476), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n944), .B(KEYINPUT108), .ZN(new_n945));
  INV_X1    g520(.A(G1996), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n752), .B(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n728), .B(G2067), .Z(new_n948));
  INV_X1    g523(.A(new_n793), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n791), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n791), .A2(new_n949), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n947), .A2(new_n948), .A3(new_n950), .A4(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(G290), .B(G1986), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n945), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT120), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n501), .A2(new_n939), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT45), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n939), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n958), .A2(new_n946), .A3(new_n943), .A4(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(G1384), .B1(new_n496), .B2(new_n500), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n943), .A2(new_n961), .ZN(new_n962));
  XOR2_X1   g537(.A(KEYINPUT58), .B(G1341), .Z(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n960), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT59), .B1(new_n965), .B2(new_n549), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT59), .ZN(new_n967));
  AOI211_X1 g542(.A(new_n967), .B(new_n548), .C1(new_n960), .C2(new_n964), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT61), .ZN(new_n970));
  XOR2_X1   g545(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n971));
  OAI21_X1  g546(.A(new_n943), .B1(new_n961), .B2(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT50), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n961), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n813), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT57), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n558), .A2(new_n565), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n536), .A2(G91), .ZN(new_n978));
  AND4_X1   g553(.A1(new_n976), .A2(new_n572), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n976), .B1(new_n566), .B2(new_n572), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(KEYINPUT56), .B(G2072), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n958), .A2(new_n943), .A3(new_n959), .A4(new_n982), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n975), .A2(new_n981), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n981), .B1(new_n975), .B2(new_n983), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n970), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n975), .A2(new_n983), .ZN(new_n987));
  INV_X1    g562(.A(new_n981), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n975), .A2(new_n981), .A3(new_n983), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(KEYINPUT61), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n969), .A2(new_n986), .A3(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT119), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n962), .A2(G2067), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n469), .A2(G40), .A3(new_n476), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(new_n956), .B2(KEYINPUT50), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n961), .A2(new_n997), .A3(new_n971), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n501), .A2(new_n939), .A3(new_n971), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(KEYINPUT111), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n996), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(G1348), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n994), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n993), .B1(new_n1003), .B2(KEYINPUT60), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1006));
  INV_X1    g581(.A(new_n994), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1006), .A2(new_n993), .A3(KEYINPUT60), .A4(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(new_n622), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1003), .A2(KEYINPUT60), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n622), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1010), .B1(new_n1011), .B2(new_n1004), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n992), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1003), .A2(new_n613), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n989), .B1(new_n1014), .B2(new_n984), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n955), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT116), .ZN(new_n1017));
  INV_X1    g592(.A(new_n971), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n956), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n961), .A2(new_n973), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT112), .B(G2090), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1019), .A2(new_n943), .A3(new_n1020), .A4(new_n1021), .ZN(new_n1022));
  AOI211_X1 g597(.A(new_n957), .B(G1384), .C1(new_n496), .C2(new_n500), .ZN(new_n1023));
  NOR3_X1   g598(.A1(new_n940), .A2(new_n1023), .A3(new_n995), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1022), .B1(new_n1024), .B2(G1971), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(G8), .ZN(new_n1026));
  XNOR2_X1  g601(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1027));
  OAI211_X1 g602(.A(G8), .B(new_n1027), .C1(new_n509), .C2(new_n520), .ZN(new_n1028));
  INV_X1    g603(.A(G8), .ZN(new_n1029));
  NOR2_X1   g604(.A1(G166), .A2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(KEYINPUT113), .A2(KEYINPUT55), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1028), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1017), .B1(new_n1026), .B2(new_n1034), .ZN(new_n1035));
  AOI211_X1 g610(.A(KEYINPUT116), .B(new_n1033), .C1(new_n1025), .C2(G8), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT109), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n1024), .B2(G1971), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n943), .B1(new_n961), .B2(new_n973), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n997), .B1(new_n961), .B2(new_n971), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(new_n998), .A3(new_n1021), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n958), .A2(new_n943), .A3(new_n959), .ZN(new_n1044));
  INV_X1    g619(.A(G1971), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1044), .A2(KEYINPUT109), .A3(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1039), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1047), .A2(G8), .A3(new_n1033), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1029), .B1(new_n943), .B2(new_n961), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n576), .A2(new_n577), .A3(G1976), .A4(new_n578), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT114), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1050), .A2(KEYINPUT114), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT52), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT52), .B1(G288), .B2(new_n772), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1049), .A2(new_n1055), .A3(new_n1051), .A4(new_n1052), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  AND2_X1   g632(.A1(new_n587), .A2(new_n588), .ZN(new_n1058));
  INV_X1    g633(.A(G1981), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1058), .B(new_n1059), .C1(new_n583), .C2(new_n585), .ZN(new_n1060));
  OAI21_X1  g635(.A(G1981), .B1(new_n586), .B2(new_n589), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT49), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1049), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(KEYINPUT115), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1062), .A2(KEYINPUT115), .A3(new_n1063), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1057), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1048), .A2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT125), .B1(new_n1037), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1029), .B1(new_n1071), .B2(new_n1022), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT116), .B1(new_n1072), .B2(new_n1033), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1026), .A2(new_n1017), .A3(new_n1034), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT125), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(new_n1076), .A3(new_n1048), .A4(new_n1068), .ZN(new_n1077));
  AND2_X1   g652(.A1(new_n1070), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n959), .A2(KEYINPUT117), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT117), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n961), .A2(new_n1080), .A3(KEYINPUT45), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1079), .A2(new_n958), .A3(new_n943), .A4(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(G1966), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n996), .A2(new_n1000), .A3(new_n732), .A4(new_n998), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1084), .A2(G168), .A3(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(G8), .ZN(new_n1087));
  AOI21_X1  g662(.A(G168), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT51), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1086), .A2(new_n1091), .A3(G8), .ZN(new_n1092));
  AND3_X1   g667(.A1(new_n1089), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1090), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1093), .A2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1096), .B1(new_n1044), .B2(G2078), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1001), .A2(new_n803), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n995), .A2(KEYINPUT123), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT123), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n469), .A2(new_n1100), .A3(G40), .A4(new_n476), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1096), .A2(G2078), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1099), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT124), .ZN(new_n1104));
  NOR4_X1   g679(.A1(new_n1103), .A2(new_n1104), .A3(new_n940), .A4(new_n1023), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1099), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n940), .A2(new_n1023), .ZN(new_n1107));
  AOI21_X1  g682(.A(KEYINPUT124), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1097), .B(new_n1098), .C1(new_n1105), .C2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G171), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT126), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1109), .A2(KEYINPUT126), .A3(G171), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n1115));
  INV_X1    g690(.A(G2078), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT53), .B1(new_n1024), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT122), .ZN(new_n1118));
  AOI21_X1  g693(.A(G1961), .B1(new_n1042), .B2(new_n998), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n995), .B1(new_n956), .B2(new_n957), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1120), .A2(new_n1079), .A3(new_n1081), .A4(new_n1102), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1118), .B1(new_n1119), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1098), .A2(KEYINPUT122), .A3(new_n1121), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1117), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1115), .B1(new_n1125), .B2(G301), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1119), .A2(new_n1117), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1127), .B(G301), .C1(new_n1108), .C2(new_n1105), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1128), .B1(new_n1125), .B2(G301), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1114), .A2(new_n1126), .B1(new_n1129), .B2(new_n1115), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1016), .A2(new_n1078), .A3(new_n1095), .A4(new_n1130), .ZN(new_n1131));
  NOR3_X1   g706(.A1(new_n1013), .A2(new_n955), .A3(new_n1015), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1134));
  NOR2_X1   g709(.A1(G288), .A2(G1976), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1134), .A2(new_n1135), .B1(new_n1059), .B2(new_n590), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1049), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1068), .ZN(new_n1138));
  OAI22_X1  g713(.A1(new_n1136), .A2(new_n1137), .B1(new_n1138), .B2(new_n1048), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1033), .B1(new_n1047), .B2(G8), .ZN(new_n1140));
  NOR2_X1   g715(.A1(G286), .A2(new_n1029), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1085), .ZN(new_n1143));
  OAI211_X1 g718(.A(KEYINPUT63), .B(new_n1141), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  NOR4_X1   g719(.A1(new_n1069), .A2(new_n1140), .A3(KEYINPUT118), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT118), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1048), .A2(new_n1068), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1047), .A2(G8), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1144), .B1(new_n1034), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1146), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT63), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1147), .A2(new_n1075), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1141), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1152), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1139), .B1(new_n1151), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1125), .A2(G301), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1070), .A2(new_n1077), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT62), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1159), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1089), .A2(new_n1092), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(KEYINPUT121), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1089), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1162), .A2(KEYINPUT62), .A3(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1158), .A2(new_n1160), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1156), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n954), .B1(new_n1133), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT46), .ZN(new_n1168));
  INV_X1    g743(.A(new_n945), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1168), .B1(new_n1169), .B2(G1996), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n945), .A2(KEYINPUT46), .A3(new_n946), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n753), .A2(new_n948), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n1170), .B(new_n1171), .C1(new_n1169), .C2(new_n1172), .ZN(new_n1173));
  XOR2_X1   g748(.A(new_n1173), .B(KEYINPUT127), .Z(new_n1174));
  XNOR2_X1  g749(.A(new_n1174), .B(KEYINPUT47), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n947), .A2(new_n948), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n1176), .A2(new_n950), .B1(G2067), .B2(new_n728), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n945), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n1169), .A2(G1986), .A3(G290), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1179), .A2(KEYINPUT48), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n952), .A2(new_n945), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NOR2_X1   g757(.A1(new_n1179), .A2(KEYINPUT48), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1178), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1175), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1167), .A2(new_n1185), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g761(.A1(G229), .A2(new_n460), .A3(G401), .A4(G227), .ZN(new_n1188));
  NAND3_X1  g762(.A1(new_n859), .A2(new_n929), .A3(new_n1188), .ZN(G225));
  INV_X1    g763(.A(G225), .ZN(G308));
endmodule


