

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U549 ( .A1(G2105), .A2(n543), .ZN(n890) );
  AND2_X1 U550 ( .A1(n766), .A2(n515), .ZN(n803) );
  BUF_X1 U551 ( .A(n561), .Z(n544) );
  NOR2_X1 U552 ( .A1(G2105), .A2(G2104), .ZN(n537) );
  NAND2_X2 U553 ( .A1(G8), .A2(n713), .ZN(n765) );
  NAND2_X2 U554 ( .A1(n769), .A2(n767), .ZN(n713) );
  NOR2_X2 U555 ( .A1(G164), .A2(G1384), .ZN(n769) );
  NOR2_X2 U556 ( .A1(n553), .A2(n552), .ZN(G164) );
  XNOR2_X1 U557 ( .A(n761), .B(KEYINPUT101), .ZN(n766) );
  NOR2_X1 U558 ( .A1(G651), .A2(G543), .ZN(n640) );
  OR2_X1 U559 ( .A1(n914), .A2(n741), .ZN(n513) );
  XOR2_X1 U560 ( .A(KEYINPUT98), .B(KEYINPUT32), .Z(n514) );
  OR2_X1 U561 ( .A1(n765), .A2(n764), .ZN(n515) );
  XNOR2_X1 U562 ( .A(n713), .B(KEYINPUT91), .ZN(n692) );
  INV_X1 U563 ( .A(n692), .ZN(n706) );
  NOR2_X1 U564 ( .A1(n717), .A2(G168), .ZN(n718) );
  NOR2_X1 U565 ( .A1(n724), .A2(n723), .ZN(n735) );
  XNOR2_X1 U566 ( .A(n733), .B(n514), .ZN(n753) );
  NOR2_X1 U567 ( .A1(n679), .A2(n678), .ZN(n767) );
  INV_X1 U568 ( .A(G651), .ZN(n520) );
  INV_X1 U569 ( .A(KEYINPUT17), .ZN(n536) );
  NOR2_X1 U570 ( .A1(G651), .A2(n616), .ZN(n646) );
  NAND2_X1 U571 ( .A1(n887), .A2(G137), .ZN(n566) );
  NAND2_X1 U572 ( .A1(n640), .A2(G89), .ZN(n516) );
  XNOR2_X1 U573 ( .A(n516), .B(KEYINPUT4), .ZN(n518) );
  XOR2_X1 U574 ( .A(KEYINPUT0), .B(G543), .Z(n616) );
  NOR2_X1 U575 ( .A1(n616), .A2(n520), .ZN(n637) );
  NAND2_X1 U576 ( .A1(G76), .A2(n637), .ZN(n517) );
  NAND2_X1 U577 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U578 ( .A(KEYINPUT5), .B(n519), .ZN(n528) );
  NAND2_X1 U579 ( .A1(n646), .A2(G51), .ZN(n524) );
  NOR2_X1 U580 ( .A1(G543), .A2(n520), .ZN(n521) );
  XOR2_X1 U581 ( .A(KEYINPUT66), .B(n521), .Z(n522) );
  XNOR2_X2 U582 ( .A(KEYINPUT1), .B(n522), .ZN(n641) );
  NAND2_X1 U583 ( .A1(G63), .A2(n641), .ZN(n523) );
  NAND2_X1 U584 ( .A1(n524), .A2(n523), .ZN(n526) );
  XOR2_X1 U585 ( .A(KEYINPUT6), .B(KEYINPUT72), .Z(n525) );
  XNOR2_X1 U586 ( .A(n526), .B(n525), .ZN(n527) );
  NAND2_X1 U587 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U588 ( .A(KEYINPUT7), .B(n529), .ZN(G168) );
  INV_X1 U589 ( .A(G2104), .ZN(n532) );
  AND2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n891) );
  NAND2_X1 U591 ( .A1(G111), .A2(n891), .ZN(n530) );
  XOR2_X1 U592 ( .A(KEYINPUT76), .B(n530), .Z(n542) );
  INV_X1 U593 ( .A(KEYINPUT64), .ZN(n531) );
  NAND2_X1 U594 ( .A1(G2104), .A2(n531), .ZN(n534) );
  NAND2_X1 U595 ( .A1(n532), .A2(KEYINPUT64), .ZN(n533) );
  NAND2_X1 U596 ( .A1(n534), .A2(n533), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n890), .A2(G123), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n535), .B(KEYINPUT18), .ZN(n539) );
  XNOR2_X2 U599 ( .A(n537), .B(n536), .ZN(n887) );
  NAND2_X1 U600 ( .A1(G135), .A2(n887), .ZN(n538) );
  NAND2_X1 U601 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U602 ( .A(KEYINPUT75), .B(n540), .Z(n541) );
  NOR2_X1 U603 ( .A1(n542), .A2(n541), .ZN(n546) );
  NOR2_X2 U604 ( .A1(G2105), .A2(n543), .ZN(n561) );
  NAND2_X1 U605 ( .A1(n544), .A2(G99), .ZN(n545) );
  NAND2_X1 U606 ( .A1(n546), .A2(n545), .ZN(n979) );
  XNOR2_X1 U607 ( .A(G2096), .B(n979), .ZN(n547) );
  OR2_X1 U608 ( .A1(G2100), .A2(n547), .ZN(G156) );
  AND2_X1 U609 ( .A1(G126), .A2(n890), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G138), .A2(n887), .ZN(n551) );
  NAND2_X1 U611 ( .A1(G114), .A2(n891), .ZN(n549) );
  NAND2_X1 U612 ( .A1(G102), .A2(n561), .ZN(n548) );
  AND2_X1 U613 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U614 ( .A1(n551), .A2(n550), .ZN(n552) );
  INV_X1 U615 ( .A(G57), .ZN(G237) );
  INV_X1 U616 ( .A(G132), .ZN(G219) );
  INV_X1 U617 ( .A(G82), .ZN(G220) );
  NAND2_X1 U618 ( .A1(n646), .A2(G52), .ZN(n555) );
  NAND2_X1 U619 ( .A1(G64), .A2(n641), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n555), .A2(n554), .ZN(n560) );
  NAND2_X1 U621 ( .A1(G77), .A2(n637), .ZN(n557) );
  NAND2_X1 U622 ( .A1(G90), .A2(n640), .ZN(n556) );
  NAND2_X1 U623 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(G171) );
  XOR2_X1 U626 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U627 ( .A1(n891), .A2(G113), .ZN(n564) );
  NAND2_X1 U628 ( .A1(G101), .A2(n561), .ZN(n562) );
  XOR2_X1 U629 ( .A(KEYINPUT23), .B(n562), .Z(n563) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n678) );
  NAND2_X1 U631 ( .A1(G125), .A2(n890), .ZN(n565) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n677) );
  NOR2_X1 U633 ( .A1(n678), .A2(n677), .ZN(G160) );
  NAND2_X1 U634 ( .A1(G94), .A2(G452), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n567), .B(KEYINPUT67), .ZN(G173) );
  NAND2_X1 U636 ( .A1(G7), .A2(G661), .ZN(n568) );
  XNOR2_X1 U637 ( .A(n568), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U638 ( .A(G223), .B(KEYINPUT68), .Z(n831) );
  NAND2_X1 U639 ( .A1(n831), .A2(G567), .ZN(n569) );
  XOR2_X1 U640 ( .A(KEYINPUT11), .B(n569), .Z(G234) );
  NAND2_X1 U641 ( .A1(G56), .A2(n641), .ZN(n570) );
  XNOR2_X1 U642 ( .A(KEYINPUT14), .B(n570), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n640), .A2(G81), .ZN(n571) );
  XNOR2_X1 U644 ( .A(n571), .B(KEYINPUT12), .ZN(n573) );
  NAND2_X1 U645 ( .A1(G68), .A2(n637), .ZN(n572) );
  NAND2_X1 U646 ( .A1(n573), .A2(n572), .ZN(n574) );
  XNOR2_X1 U647 ( .A(KEYINPUT13), .B(n574), .ZN(n575) );
  NAND2_X1 U648 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U649 ( .A(n577), .B(KEYINPUT69), .ZN(n579) );
  NAND2_X1 U650 ( .A1(n646), .A2(G43), .ZN(n578) );
  NAND2_X1 U651 ( .A1(n579), .A2(n578), .ZN(n931) );
  INV_X1 U652 ( .A(G860), .ZN(n600) );
  OR2_X1 U653 ( .A1(n931), .A2(n600), .ZN(G153) );
  INV_X1 U654 ( .A(G171), .ZN(G301) );
  NAND2_X1 U655 ( .A1(n640), .A2(G92), .ZN(n581) );
  NAND2_X1 U656 ( .A1(G66), .A2(n641), .ZN(n580) );
  NAND2_X1 U657 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U658 ( .A(KEYINPUT70), .B(n582), .ZN(n586) );
  NAND2_X1 U659 ( .A1(G79), .A2(n637), .ZN(n584) );
  NAND2_X1 U660 ( .A1(G54), .A2(n646), .ZN(n583) );
  NAND2_X1 U661 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U662 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X2 U663 ( .A(KEYINPUT15), .B(n587), .Z(n927) );
  NOR2_X1 U664 ( .A1(n927), .A2(G868), .ZN(n588) );
  XNOR2_X1 U665 ( .A(n588), .B(KEYINPUT71), .ZN(n590) );
  NAND2_X1 U666 ( .A1(G868), .A2(G301), .ZN(n589) );
  NAND2_X1 U667 ( .A1(n590), .A2(n589), .ZN(G284) );
  NAND2_X1 U668 ( .A1(n646), .A2(G53), .ZN(n592) );
  NAND2_X1 U669 ( .A1(G65), .A2(n641), .ZN(n591) );
  NAND2_X1 U670 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U671 ( .A1(G78), .A2(n637), .ZN(n594) );
  NAND2_X1 U672 ( .A1(G91), .A2(n640), .ZN(n593) );
  NAND2_X1 U673 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U674 ( .A1(n596), .A2(n595), .ZN(n915) );
  INV_X1 U675 ( .A(n915), .ZN(G299) );
  XNOR2_X1 U676 ( .A(KEYINPUT73), .B(G868), .ZN(n597) );
  NOR2_X1 U677 ( .A1(G286), .A2(n597), .ZN(n599) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U679 ( .A1(n599), .A2(n598), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n600), .A2(G559), .ZN(n601) );
  NAND2_X1 U681 ( .A1(n601), .A2(n927), .ZN(n602) );
  XNOR2_X1 U682 ( .A(n602), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U683 ( .A1(n927), .A2(G868), .ZN(n603) );
  NOR2_X1 U684 ( .A1(G559), .A2(n603), .ZN(n604) );
  XNOR2_X1 U685 ( .A(n604), .B(KEYINPUT74), .ZN(n606) );
  NOR2_X1 U686 ( .A1(n931), .A2(G868), .ZN(n605) );
  NOR2_X1 U687 ( .A1(n606), .A2(n605), .ZN(G282) );
  NAND2_X1 U688 ( .A1(n640), .A2(G93), .ZN(n608) );
  NAND2_X1 U689 ( .A1(G67), .A2(n641), .ZN(n607) );
  NAND2_X1 U690 ( .A1(n608), .A2(n607), .ZN(n611) );
  NAND2_X1 U691 ( .A1(G55), .A2(n646), .ZN(n609) );
  XNOR2_X1 U692 ( .A(KEYINPUT77), .B(n609), .ZN(n610) );
  NOR2_X1 U693 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n637), .A2(G80), .ZN(n612) );
  NAND2_X1 U695 ( .A1(n613), .A2(n612), .ZN(n659) );
  NAND2_X1 U696 ( .A1(n927), .A2(G559), .ZN(n656) );
  XNOR2_X1 U697 ( .A(n931), .B(n656), .ZN(n614) );
  NOR2_X1 U698 ( .A1(G860), .A2(n614), .ZN(n615) );
  XOR2_X1 U699 ( .A(n659), .B(n615), .Z(G145) );
  NAND2_X1 U700 ( .A1(G87), .A2(n616), .ZN(n618) );
  NAND2_X1 U701 ( .A1(G74), .A2(G651), .ZN(n617) );
  NAND2_X1 U702 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U703 ( .A1(n641), .A2(n619), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n646), .A2(G49), .ZN(n620) );
  NAND2_X1 U705 ( .A1(n621), .A2(n620), .ZN(G288) );
  NAND2_X1 U706 ( .A1(G88), .A2(n640), .ZN(n622) );
  XNOR2_X1 U707 ( .A(n622), .B(KEYINPUT80), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n641), .A2(G62), .ZN(n623) );
  XOR2_X1 U709 ( .A(KEYINPUT79), .B(n623), .Z(n624) );
  NAND2_X1 U710 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U711 ( .A1(G75), .A2(n637), .ZN(n627) );
  NAND2_X1 U712 ( .A1(G50), .A2(n646), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U714 ( .A1(n629), .A2(n628), .ZN(G166) );
  NAND2_X1 U715 ( .A1(n646), .A2(G47), .ZN(n631) );
  NAND2_X1 U716 ( .A1(G60), .A2(n641), .ZN(n630) );
  NAND2_X1 U717 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U718 ( .A1(G72), .A2(n637), .ZN(n632) );
  XNOR2_X1 U719 ( .A(KEYINPUT65), .B(n632), .ZN(n633) );
  NOR2_X1 U720 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U721 ( .A1(n640), .A2(G85), .ZN(n635) );
  NAND2_X1 U722 ( .A1(n636), .A2(n635), .ZN(G290) );
  XOR2_X1 U723 ( .A(KEYINPUT78), .B(KEYINPUT2), .Z(n639) );
  NAND2_X1 U724 ( .A1(G73), .A2(n637), .ZN(n638) );
  XNOR2_X1 U725 ( .A(n639), .B(n638), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n640), .A2(G86), .ZN(n643) );
  NAND2_X1 U727 ( .A1(G61), .A2(n641), .ZN(n642) );
  NAND2_X1 U728 ( .A1(n643), .A2(n642), .ZN(n644) );
  NOR2_X1 U729 ( .A1(n645), .A2(n644), .ZN(n648) );
  NAND2_X1 U730 ( .A1(n646), .A2(G48), .ZN(n647) );
  NAND2_X1 U731 ( .A1(n648), .A2(n647), .ZN(G305) );
  XNOR2_X1 U732 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n650) );
  XNOR2_X1 U733 ( .A(G288), .B(G166), .ZN(n649) );
  XNOR2_X1 U734 ( .A(n650), .B(n649), .ZN(n653) );
  XOR2_X1 U735 ( .A(G290), .B(n931), .Z(n651) );
  XNOR2_X1 U736 ( .A(n659), .B(n651), .ZN(n652) );
  XNOR2_X1 U737 ( .A(n653), .B(n652), .ZN(n655) );
  XNOR2_X1 U738 ( .A(G305), .B(n915), .ZN(n654) );
  XNOR2_X1 U739 ( .A(n655), .B(n654), .ZN(n902) );
  XOR2_X1 U740 ( .A(n902), .B(n656), .Z(n657) );
  NAND2_X1 U741 ( .A1(G868), .A2(n657), .ZN(n661) );
  INV_X1 U742 ( .A(G868), .ZN(n658) );
  NAND2_X1 U743 ( .A1(n659), .A2(n658), .ZN(n660) );
  NAND2_X1 U744 ( .A1(n661), .A2(n660), .ZN(G295) );
  NAND2_X1 U745 ( .A1(G2078), .A2(G2084), .ZN(n662) );
  XOR2_X1 U746 ( .A(KEYINPUT20), .B(n662), .Z(n663) );
  NAND2_X1 U747 ( .A1(G2090), .A2(n663), .ZN(n664) );
  XNOR2_X1 U748 ( .A(KEYINPUT21), .B(n664), .ZN(n665) );
  NAND2_X1 U749 ( .A1(n665), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U750 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U751 ( .A1(G220), .A2(G219), .ZN(n666) );
  XOR2_X1 U752 ( .A(KEYINPUT22), .B(n666), .Z(n667) );
  NOR2_X1 U753 ( .A1(G218), .A2(n667), .ZN(n668) );
  NAND2_X1 U754 ( .A1(G96), .A2(n668), .ZN(n911) );
  NAND2_X1 U755 ( .A1(G2106), .A2(n911), .ZN(n672) );
  NAND2_X1 U756 ( .A1(G69), .A2(G120), .ZN(n669) );
  NOR2_X1 U757 ( .A1(G237), .A2(n669), .ZN(n670) );
  NAND2_X1 U758 ( .A1(G108), .A2(n670), .ZN(n912) );
  NAND2_X1 U759 ( .A1(G567), .A2(n912), .ZN(n671) );
  NAND2_X1 U760 ( .A1(n672), .A2(n671), .ZN(n837) );
  NAND2_X1 U761 ( .A1(G483), .A2(G661), .ZN(n673) );
  NOR2_X1 U762 ( .A1(n837), .A2(n673), .ZN(n835) );
  NAND2_X1 U763 ( .A1(G36), .A2(n835), .ZN(n674) );
  XNOR2_X1 U764 ( .A(n674), .B(KEYINPUT82), .ZN(G176) );
  INV_X1 U765 ( .A(G166), .ZN(G303) );
  INV_X1 U766 ( .A(G40), .ZN(n676) );
  OR2_X1 U767 ( .A1(n677), .A2(n676), .ZN(n679) );
  NAND2_X1 U768 ( .A1(n692), .A2(G2072), .ZN(n680) );
  XNOR2_X1 U769 ( .A(n680), .B(KEYINPUT27), .ZN(n682) );
  AND2_X1 U770 ( .A1(G1956), .A2(n706), .ZN(n681) );
  NOR2_X1 U771 ( .A1(n682), .A2(n681), .ZN(n685) );
  NOR2_X1 U772 ( .A1(n685), .A2(n915), .ZN(n684) );
  INV_X1 U773 ( .A(KEYINPUT28), .ZN(n683) );
  XNOR2_X1 U774 ( .A(n684), .B(n683), .ZN(n702) );
  NAND2_X1 U775 ( .A1(n915), .A2(n685), .ZN(n700) );
  INV_X1 U776 ( .A(n713), .ZN(n705) );
  AND2_X1 U777 ( .A1(n705), .A2(G1996), .ZN(n687) );
  XOR2_X1 U778 ( .A(KEYINPUT26), .B(KEYINPUT94), .Z(n686) );
  XNOR2_X1 U779 ( .A(n687), .B(n686), .ZN(n689) );
  NAND2_X1 U780 ( .A1(n713), .A2(G1341), .ZN(n688) );
  NAND2_X1 U781 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U782 ( .A1(n931), .A2(n690), .ZN(n691) );
  OR2_X1 U783 ( .A1(n927), .A2(n691), .ZN(n698) );
  NAND2_X1 U784 ( .A1(n927), .A2(n691), .ZN(n696) );
  NAND2_X1 U785 ( .A1(G2067), .A2(n692), .ZN(n694) );
  NAND2_X1 U786 ( .A1(G1348), .A2(n713), .ZN(n693) );
  NAND2_X1 U787 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U788 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U789 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U790 ( .A1(n700), .A2(n699), .ZN(n701) );
  AND2_X1 U791 ( .A1(n702), .A2(n701), .ZN(n704) );
  XNOR2_X1 U792 ( .A(KEYINPUT29), .B(KEYINPUT95), .ZN(n703) );
  XNOR2_X1 U793 ( .A(n704), .B(n703), .ZN(n712) );
  NOR2_X1 U794 ( .A1(n705), .A2(G1961), .ZN(n708) );
  XOR2_X1 U795 ( .A(G2078), .B(KEYINPUT25), .Z(n949) );
  NOR2_X1 U796 ( .A1(n949), .A2(n706), .ZN(n707) );
  NOR2_X1 U797 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U798 ( .A(n709), .B(KEYINPUT92), .ZN(n719) );
  NOR2_X1 U799 ( .A1(G301), .A2(n719), .ZN(n710) );
  XOR2_X1 U800 ( .A(KEYINPUT93), .B(n710), .Z(n711) );
  NOR2_X1 U801 ( .A1(n712), .A2(n711), .ZN(n724) );
  NOR2_X1 U802 ( .A1(G2084), .A2(n713), .ZN(n734) );
  NOR2_X1 U803 ( .A1(G1966), .A2(n765), .ZN(n736) );
  NOR2_X1 U804 ( .A1(n734), .A2(n736), .ZN(n714) );
  XNOR2_X1 U805 ( .A(n714), .B(KEYINPUT96), .ZN(n715) );
  NAND2_X1 U806 ( .A1(n715), .A2(G8), .ZN(n716) );
  XNOR2_X1 U807 ( .A(n716), .B(KEYINPUT30), .ZN(n717) );
  XNOR2_X1 U808 ( .A(n718), .B(KEYINPUT97), .ZN(n721) );
  NAND2_X1 U809 ( .A1(n719), .A2(G301), .ZN(n720) );
  AND2_X1 U810 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U811 ( .A(n722), .B(KEYINPUT31), .ZN(n723) );
  INV_X1 U812 ( .A(n735), .ZN(n725) );
  NAND2_X1 U813 ( .A1(n725), .A2(G286), .ZN(n732) );
  INV_X1 U814 ( .A(G8), .ZN(n730) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n765), .ZN(n727) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n713), .ZN(n726) );
  NOR2_X1 U817 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U818 ( .A1(G303), .A2(n728), .ZN(n729) );
  OR2_X1 U819 ( .A1(n730), .A2(n729), .ZN(n731) );
  NAND2_X1 U820 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U821 ( .A1(n734), .A2(G8), .ZN(n738) );
  NOR2_X1 U822 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U823 ( .A1(n738), .A2(n737), .ZN(n754) );
  NAND2_X1 U824 ( .A1(G1976), .A2(G288), .ZN(n740) );
  AND2_X1 U825 ( .A1(n754), .A2(n740), .ZN(n739) );
  NAND2_X1 U826 ( .A1(n753), .A2(n739), .ZN(n742) );
  INV_X1 U827 ( .A(n740), .ZN(n914) );
  NOR2_X1 U828 ( .A1(G1971), .A2(G303), .ZN(n913) );
  NOR2_X1 U829 ( .A1(G1976), .A2(G288), .ZN(n918) );
  NOR2_X1 U830 ( .A1(n913), .A2(n918), .ZN(n741) );
  AND2_X1 U831 ( .A1(n742), .A2(n513), .ZN(n743) );
  XNOR2_X1 U832 ( .A(n743), .B(KEYINPUT99), .ZN(n746) );
  INV_X1 U833 ( .A(KEYINPUT33), .ZN(n744) );
  INV_X1 U834 ( .A(n765), .ZN(n747) );
  AND2_X1 U835 ( .A1(n744), .A2(n747), .ZN(n745) );
  NAND2_X1 U836 ( .A1(n746), .A2(n745), .ZN(n750) );
  NAND2_X1 U837 ( .A1(n918), .A2(n747), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n748), .A2(KEYINPUT33), .ZN(n749) );
  NAND2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U840 ( .A(n751), .B(KEYINPUT100), .ZN(n752) );
  XOR2_X1 U841 ( .A(G1981), .B(G305), .Z(n932) );
  NAND2_X1 U842 ( .A1(n752), .A2(n932), .ZN(n760) );
  NAND2_X1 U843 ( .A1(n754), .A2(n753), .ZN(n757) );
  NOR2_X1 U844 ( .A1(G2090), .A2(G303), .ZN(n755) );
  NAND2_X1 U845 ( .A1(G8), .A2(n755), .ZN(n756) );
  NAND2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U847 ( .A1(n758), .A2(n765), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U849 ( .A1(G1981), .A2(G305), .ZN(n762) );
  XOR2_X1 U850 ( .A(n762), .B(KEYINPUT90), .Z(n763) );
  XNOR2_X1 U851 ( .A(KEYINPUT24), .B(n763), .ZN(n764) );
  INV_X1 U852 ( .A(n767), .ZN(n768) );
  NOR2_X1 U853 ( .A1(n769), .A2(n768), .ZN(n816) );
  NAND2_X1 U854 ( .A1(G140), .A2(n887), .ZN(n771) );
  NAND2_X1 U855 ( .A1(G104), .A2(n544), .ZN(n770) );
  NAND2_X1 U856 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U857 ( .A(KEYINPUT34), .B(n772), .ZN(n778) );
  NAND2_X1 U858 ( .A1(G128), .A2(n890), .ZN(n774) );
  NAND2_X1 U859 ( .A1(G116), .A2(n891), .ZN(n773) );
  NAND2_X1 U860 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U861 ( .A(KEYINPUT35), .B(n775), .Z(n776) );
  XNOR2_X1 U862 ( .A(KEYINPUT84), .B(n776), .ZN(n777) );
  NOR2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U864 ( .A(KEYINPUT36), .B(n779), .ZN(n867) );
  XOR2_X1 U865 ( .A(G2067), .B(KEYINPUT37), .Z(n780) );
  XNOR2_X1 U866 ( .A(KEYINPUT83), .B(n780), .ZN(n814) );
  NOR2_X1 U867 ( .A1(n867), .A2(n814), .ZN(n978) );
  NAND2_X1 U868 ( .A1(n816), .A2(n978), .ZN(n812) );
  NAND2_X1 U869 ( .A1(G105), .A2(n544), .ZN(n781) );
  XNOR2_X1 U870 ( .A(n781), .B(KEYINPUT38), .ZN(n782) );
  XNOR2_X1 U871 ( .A(n782), .B(KEYINPUT86), .ZN(n784) );
  NAND2_X1 U872 ( .A1(G117), .A2(n891), .ZN(n783) );
  NAND2_X1 U873 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U874 ( .A1(G141), .A2(n887), .ZN(n785) );
  XNOR2_X1 U875 ( .A(KEYINPUT87), .B(n785), .ZN(n786) );
  NOR2_X1 U876 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U877 ( .A1(G129), .A2(n890), .ZN(n788) );
  XOR2_X1 U878 ( .A(KEYINPUT85), .B(n788), .Z(n789) );
  NAND2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n871) );
  AND2_X1 U880 ( .A1(n871), .A2(G1996), .ZN(n798) );
  NAND2_X1 U881 ( .A1(G131), .A2(n887), .ZN(n792) );
  NAND2_X1 U882 ( .A1(G95), .A2(n544), .ZN(n791) );
  NAND2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U884 ( .A1(G119), .A2(n890), .ZN(n794) );
  NAND2_X1 U885 ( .A1(G107), .A2(n891), .ZN(n793) );
  NAND2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n795) );
  OR2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n884) );
  AND2_X1 U888 ( .A1(n884), .A2(G1991), .ZN(n797) );
  NOR2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n976) );
  XOR2_X1 U890 ( .A(n816), .B(KEYINPUT88), .Z(n799) );
  NOR2_X1 U891 ( .A1(n976), .A2(n799), .ZN(n808) );
  INV_X1 U892 ( .A(n808), .ZN(n800) );
  NAND2_X1 U893 ( .A1(n812), .A2(n800), .ZN(n801) );
  XOR2_X1 U894 ( .A(KEYINPUT89), .B(n801), .Z(n802) );
  NOR2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n805) );
  XNOR2_X1 U896 ( .A(G1986), .B(G290), .ZN(n920) );
  NAND2_X1 U897 ( .A1(n920), .A2(n816), .ZN(n804) );
  NAND2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n819) );
  NOR2_X1 U899 ( .A1(G1996), .A2(n871), .ZN(n982) );
  NOR2_X1 U900 ( .A1(G1991), .A2(n884), .ZN(n974) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U902 ( .A1(n974), .A2(n806), .ZN(n807) );
  NOR2_X1 U903 ( .A1(n808), .A2(n807), .ZN(n809) );
  XNOR2_X1 U904 ( .A(n809), .B(KEYINPUT102), .ZN(n810) );
  NOR2_X1 U905 ( .A1(n982), .A2(n810), .ZN(n811) );
  XNOR2_X1 U906 ( .A(KEYINPUT39), .B(n811), .ZN(n813) );
  NAND2_X1 U907 ( .A1(n813), .A2(n812), .ZN(n815) );
  NAND2_X1 U908 ( .A1(n867), .A2(n814), .ZN(n980) );
  NAND2_X1 U909 ( .A1(n815), .A2(n980), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U911 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U912 ( .A(n820), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U913 ( .A(G2454), .B(G2430), .Z(n822) );
  XNOR2_X1 U914 ( .A(G2451), .B(G2446), .ZN(n821) );
  XNOR2_X1 U915 ( .A(n822), .B(n821), .ZN(n829) );
  XOR2_X1 U916 ( .A(G2443), .B(G2427), .Z(n824) );
  XNOR2_X1 U917 ( .A(G2438), .B(KEYINPUT103), .ZN(n823) );
  XNOR2_X1 U918 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U919 ( .A(n825), .B(G2435), .Z(n827) );
  XNOR2_X1 U920 ( .A(G1341), .B(G1348), .ZN(n826) );
  XNOR2_X1 U921 ( .A(n827), .B(n826), .ZN(n828) );
  XNOR2_X1 U922 ( .A(n829), .B(n828), .ZN(n830) );
  NAND2_X1 U923 ( .A1(n830), .A2(G14), .ZN(n905) );
  XOR2_X1 U924 ( .A(KEYINPUT104), .B(n905), .Z(G401) );
  NAND2_X1 U925 ( .A1(n831), .A2(G2106), .ZN(n832) );
  XOR2_X1 U926 ( .A(KEYINPUT105), .B(n832), .Z(G217) );
  AND2_X1 U927 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U928 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n834) );
  XNOR2_X1 U930 ( .A(KEYINPUT106), .B(n834), .ZN(n836) );
  NAND2_X1 U931 ( .A1(n836), .A2(n835), .ZN(G188) );
  XNOR2_X1 U932 ( .A(KEYINPUT107), .B(n837), .ZN(G319) );
  XOR2_X1 U933 ( .A(KEYINPUT41), .B(G1966), .Z(n839) );
  XNOR2_X1 U934 ( .A(G1981), .B(G1961), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U936 ( .A(n840), .B(G2474), .Z(n842) );
  XNOR2_X1 U937 ( .A(G1996), .B(G1991), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U939 ( .A(G1956), .B(G1971), .Z(n844) );
  XNOR2_X1 U940 ( .A(G1986), .B(G1976), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n845) );
  XOR2_X1 U942 ( .A(n846), .B(n845), .Z(n848) );
  XNOR2_X1 U943 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n847) );
  XNOR2_X1 U944 ( .A(n848), .B(n847), .ZN(G229) );
  XOR2_X1 U945 ( .A(G2096), .B(G2678), .Z(n850) );
  XNOR2_X1 U946 ( .A(G2090), .B(KEYINPUT43), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U948 ( .A(n851), .B(KEYINPUT42), .Z(n853) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U950 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U951 ( .A(KEYINPUT108), .B(G2100), .Z(n855) );
  XNOR2_X1 U952 ( .A(G2078), .B(G2084), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(G227) );
  NAND2_X1 U955 ( .A1(G112), .A2(n891), .ZN(n859) );
  NAND2_X1 U956 ( .A1(G100), .A2(n544), .ZN(n858) );
  NAND2_X1 U957 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U958 ( .A(KEYINPUT112), .B(n860), .ZN(n866) );
  NAND2_X1 U959 ( .A1(G124), .A2(n890), .ZN(n861) );
  XOR2_X1 U960 ( .A(KEYINPUT111), .B(n861), .Z(n862) );
  XNOR2_X1 U961 ( .A(n862), .B(KEYINPUT44), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G136), .A2(n887), .ZN(n863) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U964 ( .A1(n866), .A2(n865), .ZN(G162) );
  XNOR2_X1 U965 ( .A(KEYINPUT48), .B(KEYINPUT114), .ZN(n869) );
  XNOR2_X1 U966 ( .A(n867), .B(KEYINPUT46), .ZN(n868) );
  XNOR2_X1 U967 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U968 ( .A(n979), .B(n870), .ZN(n873) );
  XOR2_X1 U969 ( .A(G164), .B(n871), .Z(n872) );
  XNOR2_X1 U970 ( .A(n873), .B(n872), .ZN(n883) );
  NAND2_X1 U971 ( .A1(G142), .A2(n887), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G106), .A2(n544), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U974 ( .A(n876), .B(KEYINPUT45), .ZN(n878) );
  NAND2_X1 U975 ( .A1(G118), .A2(n891), .ZN(n877) );
  NAND2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n881) );
  NAND2_X1 U977 ( .A1(G130), .A2(n890), .ZN(n879) );
  XNOR2_X1 U978 ( .A(KEYINPUT113), .B(n879), .ZN(n880) );
  NOR2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U980 ( .A(n883), .B(n882), .Z(n886) );
  XOR2_X1 U981 ( .A(G160), .B(n884), .Z(n885) );
  XNOR2_X1 U982 ( .A(n886), .B(n885), .ZN(n898) );
  NAND2_X1 U983 ( .A1(G139), .A2(n887), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G103), .A2(n544), .ZN(n888) );
  NAND2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n896) );
  NAND2_X1 U986 ( .A1(G127), .A2(n890), .ZN(n893) );
  NAND2_X1 U987 ( .A1(G115), .A2(n891), .ZN(n892) );
  NAND2_X1 U988 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U989 ( .A(KEYINPUT47), .B(n894), .Z(n895) );
  NOR2_X1 U990 ( .A1(n896), .A2(n895), .ZN(n968) );
  XNOR2_X1 U991 ( .A(G162), .B(n968), .ZN(n897) );
  XNOR2_X1 U992 ( .A(n898), .B(n897), .ZN(n899) );
  NOR2_X1 U993 ( .A1(G37), .A2(n899), .ZN(G395) );
  XOR2_X1 U994 ( .A(KEYINPUT115), .B(G171), .Z(n901) );
  XNOR2_X1 U995 ( .A(G286), .B(n927), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n903) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U998 ( .A1(G37), .A2(n904), .ZN(G397) );
  NAND2_X1 U999 ( .A1(G319), .A2(n905), .ZN(n908) );
  NOR2_X1 U1000 ( .A1(G229), .A2(G227), .ZN(n906) );
  XNOR2_X1 U1001 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1002 ( .A1(n908), .A2(n907), .ZN(n910) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n909) );
  NAND2_X1 U1004 ( .A1(n910), .A2(n909), .ZN(G225) );
  XOR2_X1 U1005 ( .A(KEYINPUT116), .B(G225), .Z(G308) );
  INV_X1 U1007 ( .A(G120), .ZN(G236) );
  INV_X1 U1008 ( .A(G96), .ZN(G221) );
  INV_X1 U1009 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1010 ( .A1(n912), .A2(n911), .ZN(G325) );
  INV_X1 U1011 ( .A(G325), .ZN(G261) );
  INV_X1 U1012 ( .A(G108), .ZN(G238) );
  NOR2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n926) );
  XNOR2_X1 U1014 ( .A(G1956), .B(n915), .ZN(n917) );
  NAND2_X1 U1015 ( .A1(G1971), .A2(G303), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n924) );
  XNOR2_X1 U1017 ( .A(G171), .B(G1961), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(KEYINPUT122), .B(n918), .ZN(n919) );
  NOR2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n921) );
  NAND2_X1 U1020 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1021 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n930) );
  INV_X1 U1023 ( .A(n927), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(G1348), .B(n928), .ZN(n929) );
  NOR2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n939) );
  XNOR2_X1 U1026 ( .A(n931), .B(G1341), .ZN(n937) );
  XNOR2_X1 U1027 ( .A(G168), .B(G1966), .ZN(n933) );
  NAND2_X1 U1028 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1029 ( .A(n934), .B(KEYINPUT121), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(KEYINPUT57), .B(n935), .ZN(n936) );
  NOR2_X1 U1031 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n942) );
  XNOR2_X1 U1033 ( .A(G16), .B(KEYINPUT120), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(n940), .B(KEYINPUT56), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1036 ( .A(n943), .B(KEYINPUT123), .ZN(n967) );
  INV_X1 U1037 ( .A(KEYINPUT55), .ZN(n991) );
  XNOR2_X1 U1038 ( .A(G2084), .B(G34), .ZN(n944) );
  XNOR2_X1 U1039 ( .A(n944), .B(KEYINPUT54), .ZN(n958) );
  XOR2_X1 U1040 ( .A(G2072), .B(G33), .Z(n945) );
  NAND2_X1 U1041 ( .A1(n945), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1042 ( .A(G32), .B(G1996), .ZN(n946) );
  XNOR2_X1 U1043 ( .A(n946), .B(KEYINPUT119), .ZN(n953) );
  XOR2_X1 U1044 ( .A(G2067), .B(G26), .Z(n948) );
  XOR2_X1 U1045 ( .A(G1991), .B(G25), .Z(n947) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(G27), .B(n949), .ZN(n950) );
  NOR2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1049 ( .A1(n953), .A2(n952), .ZN(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(n956), .B(KEYINPUT53), .ZN(n957) );
  NOR2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1053 ( .A(G2090), .B(KEYINPUT118), .Z(n959) );
  XNOR2_X1 U1054 ( .A(G35), .B(n959), .ZN(n960) );
  NAND2_X1 U1055 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1056 ( .A(n991), .B(n962), .ZN(n964) );
  INV_X1 U1057 ( .A(G29), .ZN(n963) );
  NAND2_X1 U1058 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n965), .ZN(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n995) );
  XNOR2_X1 U1061 ( .A(G164), .B(G2078), .ZN(n971) );
  XOR2_X1 U1062 ( .A(G2072), .B(n968), .Z(n969) );
  XNOR2_X1 U1063 ( .A(KEYINPUT117), .B(n969), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n972), .B(KEYINPUT50), .ZN(n989) );
  XOR2_X1 U1066 ( .A(G160), .B(G2084), .Z(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n987) );
  NAND2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n985) );
  XOR2_X1 U1071 ( .A(G2090), .B(G162), .Z(n981) );
  NOR2_X1 U1072 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1073 ( .A(n983), .B(KEYINPUT51), .ZN(n984) );
  NOR2_X1 U1074 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1075 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(KEYINPUT52), .B(n990), .ZN(n992) );
  NAND2_X1 U1078 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1079 ( .A1(n993), .A2(G29), .ZN(n994) );
  NAND2_X1 U1080 ( .A1(n995), .A2(n994), .ZN(n1022) );
  XOR2_X1 U1081 ( .A(G1961), .B(G5), .Z(n1006) );
  XNOR2_X1 U1082 ( .A(G1348), .B(KEYINPUT59), .ZN(n996) );
  XNOR2_X1 U1083 ( .A(n996), .B(G4), .ZN(n1000) );
  XNOR2_X1 U1084 ( .A(G1341), .B(G19), .ZN(n998) );
  XNOR2_X1 U1085 ( .A(G1956), .B(G20), .ZN(n997) );
  NOR2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1003) );
  XNOR2_X1 U1088 ( .A(KEYINPUT124), .B(G1981), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(G6), .B(n1001), .ZN(n1002) );
  NOR2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XNOR2_X1 U1091 ( .A(KEYINPUT60), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1092 ( .A1(n1006), .A2(n1005), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(G21), .B(G1966), .ZN(n1007) );
  NOR2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1095 ( .A(KEYINPUT125), .B(n1009), .Z(n1017) );
  XOR2_X1 U1096 ( .A(G1971), .B(G22), .Z(n1012) );
  XOR2_X1 U1097 ( .A(G23), .B(KEYINPUT126), .Z(n1010) );
  XNOR2_X1 U1098 ( .A(n1010), .B(G1976), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1100 ( .A(G24), .B(G1986), .ZN(n1013) );
  NOR2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(KEYINPUT58), .B(n1015), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XOR2_X1 U1104 ( .A(n1018), .B(KEYINPUT61), .Z(n1019) );
  XNOR2_X1 U1105 ( .A(KEYINPUT127), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1106 ( .A1(G16), .A2(n1020), .ZN(n1021) );
  NOR2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(n1023), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

