

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592;

  XNOR2_X1 U326 ( .A(n359), .B(n339), .ZN(n340) );
  XNOR2_X1 U327 ( .A(n405), .B(n404), .ZN(n406) );
  NOR2_X1 U328 ( .A1(n370), .A2(n369), .ZN(n371) );
  XNOR2_X1 U329 ( .A(n343), .B(n342), .ZN(n472) );
  XNOR2_X1 U330 ( .A(n438), .B(n294), .ZN(n342) );
  XNOR2_X1 U331 ( .A(n407), .B(n406), .ZN(n415) );
  XOR2_X1 U332 ( .A(n363), .B(n362), .Z(n541) );
  XNOR2_X1 U333 ( .A(n486), .B(KEYINPUT38), .ZN(n516) );
  XOR2_X1 U334 ( .A(n331), .B(n330), .Z(n532) );
  AND2_X1 U335 ( .A1(G226GAT), .A2(G233GAT), .ZN(n294) );
  XOR2_X1 U336 ( .A(n423), .B(n422), .Z(n295) );
  XOR2_X1 U337 ( .A(G155GAT), .B(KEYINPUT2), .Z(n296) );
  XOR2_X1 U338 ( .A(n302), .B(G106GAT), .Z(n297) );
  XOR2_X1 U339 ( .A(G64GAT), .B(KEYINPUT74), .Z(n298) );
  XNOR2_X1 U340 ( .A(KEYINPUT45), .B(KEYINPUT66), .ZN(n456) );
  AND2_X1 U341 ( .A1(n467), .A2(n466), .ZN(n468) );
  INV_X1 U342 ( .A(n426), .ZN(n413) );
  XNOR2_X1 U343 ( .A(n407), .B(n338), .ZN(n339) );
  XNOR2_X1 U344 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U345 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U346 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U347 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U348 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U349 ( .A(n311), .B(n310), .ZN(n476) );
  XOR2_X1 U350 ( .A(n417), .B(n416), .Z(n566) );
  XNOR2_X1 U351 ( .A(KEYINPUT41), .B(n583), .ZN(n557) );
  NOR2_X1 U352 ( .A1(n485), .A2(n503), .ZN(n486) );
  INV_X1 U353 ( .A(G43GAT), .ZN(n491) );
  INV_X1 U354 ( .A(G29GAT), .ZN(n487) );
  XNOR2_X1 U355 ( .A(n495), .B(KEYINPUT122), .ZN(n496) );
  XNOR2_X1 U356 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n452) );
  XNOR2_X1 U357 ( .A(G92GAT), .B(KEYINPUT112), .ZN(n454) );
  XNOR2_X1 U358 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U359 ( .A(n497), .B(n496), .ZN(G1350GAT) );
  XNOR2_X1 U360 ( .A(n455), .B(n454), .ZN(G1337GAT) );
  XNOR2_X1 U361 ( .A(KEYINPUT3), .B(KEYINPUT89), .ZN(n299) );
  XNOR2_X1 U362 ( .A(n296), .B(n299), .ZN(n323) );
  XOR2_X1 U363 ( .A(KEYINPUT22), .B(n323), .Z(n301) );
  NAND2_X1 U364 ( .A1(G228GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U365 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U366 ( .A(G141GAT), .B(G22GAT), .Z(n439) );
  XNOR2_X1 U367 ( .A(n439), .B(G218GAT), .ZN(n303) );
  XNOR2_X1 U368 ( .A(n297), .B(n303), .ZN(n305) );
  XNOR2_X1 U369 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n304) );
  XNOR2_X1 U370 ( .A(n304), .B(G211GAT), .ZN(n333) );
  XOR2_X1 U371 ( .A(n305), .B(n333), .Z(n311) );
  XOR2_X1 U372 ( .A(G50GAT), .B(G162GAT), .Z(n411) );
  XOR2_X1 U373 ( .A(G148GAT), .B(G78GAT), .Z(n428) );
  XNOR2_X1 U374 ( .A(n411), .B(n428), .ZN(n309) );
  XOR2_X1 U375 ( .A(KEYINPUT23), .B(G204GAT), .Z(n307) );
  XNOR2_X1 U376 ( .A(KEYINPUT24), .B(KEYINPUT90), .ZN(n306) );
  XNOR2_X1 U377 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U378 ( .A(KEYINPUT28), .B(n476), .ZN(n375) );
  INV_X1 U379 ( .A(n375), .ZN(n527) );
  XOR2_X1 U380 ( .A(KEYINPUT1), .B(KEYINPUT91), .Z(n313) );
  XNOR2_X1 U381 ( .A(G1GAT), .B(KEYINPUT92), .ZN(n312) );
  XNOR2_X1 U382 ( .A(n313), .B(n312), .ZN(n331) );
  XOR2_X1 U383 ( .A(G85GAT), .B(G148GAT), .Z(n315) );
  XNOR2_X1 U384 ( .A(G127GAT), .B(G120GAT), .ZN(n314) );
  XNOR2_X1 U385 ( .A(n315), .B(n314), .ZN(n319) );
  XOR2_X1 U386 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n317) );
  XNOR2_X1 U387 ( .A(G141GAT), .B(KEYINPUT5), .ZN(n316) );
  XNOR2_X1 U388 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U389 ( .A(n319), .B(n318), .Z(n329) );
  XNOR2_X1 U390 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n320) );
  XNOR2_X1 U391 ( .A(n320), .B(KEYINPUT81), .ZN(n344) );
  XOR2_X1 U392 ( .A(n344), .B(G57GAT), .Z(n322) );
  NAND2_X1 U393 ( .A1(G225GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U394 ( .A(n322), .B(n321), .ZN(n327) );
  XOR2_X1 U395 ( .A(G134GAT), .B(KEYINPUT76), .Z(n410) );
  XOR2_X1 U396 ( .A(n410), .B(G162GAT), .Z(n325) );
  XNOR2_X1 U397 ( .A(G29GAT), .B(n323), .ZN(n324) );
  XNOR2_X1 U398 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U399 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U400 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U401 ( .A(G176GAT), .B(G204GAT), .ZN(n332) );
  XNOR2_X1 U402 ( .A(n298), .B(n332), .ZN(n423) );
  XNOR2_X1 U403 ( .A(n333), .B(n423), .ZN(n341) );
  XOR2_X1 U404 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n335) );
  XNOR2_X1 U405 ( .A(KEYINPUT88), .B(G183GAT), .ZN(n334) );
  XNOR2_X1 U406 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U407 ( .A(KEYINPUT19), .B(n336), .Z(n359) );
  XNOR2_X1 U408 ( .A(G36GAT), .B(G190GAT), .ZN(n337) );
  XNOR2_X1 U409 ( .A(n337), .B(G218GAT), .ZN(n407) );
  XOR2_X1 U410 ( .A(KEYINPUT93), .B(G92GAT), .Z(n338) );
  XNOR2_X1 U411 ( .A(n341), .B(n340), .ZN(n343) );
  XOR2_X1 U412 ( .A(G169GAT), .B(G8GAT), .Z(n438) );
  INV_X1 U413 ( .A(n472), .ZN(n523) );
  XOR2_X1 U414 ( .A(G15GAT), .B(G127GAT), .Z(n382) );
  XOR2_X1 U415 ( .A(n382), .B(n344), .Z(n346) );
  NAND2_X1 U416 ( .A1(G227GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U417 ( .A(n346), .B(n345), .ZN(n363) );
  XOR2_X1 U418 ( .A(KEYINPUT84), .B(KEYINPUT20), .Z(n348) );
  XNOR2_X1 U419 ( .A(G169GAT), .B(KEYINPUT85), .ZN(n347) );
  XNOR2_X1 U420 ( .A(n348), .B(n347), .ZN(n352) );
  XOR2_X1 U421 ( .A(G176GAT), .B(KEYINPUT64), .Z(n350) );
  XNOR2_X1 U422 ( .A(KEYINPUT83), .B(KEYINPUT87), .ZN(n349) );
  XNOR2_X1 U423 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U424 ( .A(n352), .B(n351), .Z(n361) );
  XOR2_X1 U425 ( .A(KEYINPUT86), .B(KEYINPUT82), .Z(n354) );
  XNOR2_X1 U426 ( .A(G134GAT), .B(G99GAT), .ZN(n353) );
  XNOR2_X1 U427 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U428 ( .A(n355), .B(G190GAT), .Z(n357) );
  XOR2_X1 U429 ( .A(G120GAT), .B(G71GAT), .Z(n422) );
  XNOR2_X1 U430 ( .A(G43GAT), .B(n422), .ZN(n356) );
  XNOR2_X1 U431 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U432 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U433 ( .A(n361), .B(n360), .ZN(n362) );
  NAND2_X1 U434 ( .A1(n523), .A2(n541), .ZN(n364) );
  NAND2_X1 U435 ( .A1(n364), .A2(n476), .ZN(n365) );
  XNOR2_X1 U436 ( .A(n365), .B(KEYINPUT25), .ZN(n366) );
  XNOR2_X1 U437 ( .A(n366), .B(KEYINPUT98), .ZN(n370) );
  XNOR2_X1 U438 ( .A(n523), .B(KEYINPUT27), .ZN(n373) );
  NOR2_X1 U439 ( .A1(n541), .A2(n476), .ZN(n368) );
  XNOR2_X1 U440 ( .A(KEYINPUT26), .B(KEYINPUT97), .ZN(n367) );
  XOR2_X1 U441 ( .A(n368), .B(n367), .Z(n576) );
  AND2_X1 U442 ( .A1(n373), .A2(n576), .ZN(n369) );
  XOR2_X1 U443 ( .A(KEYINPUT99), .B(n371), .Z(n372) );
  NOR2_X1 U444 ( .A1(n532), .A2(n372), .ZN(n379) );
  NAND2_X1 U445 ( .A1(n373), .A2(n532), .ZN(n374) );
  XOR2_X1 U446 ( .A(KEYINPUT94), .B(n374), .Z(n553) );
  NAND2_X1 U447 ( .A1(n375), .A2(n553), .ZN(n539) );
  XOR2_X1 U448 ( .A(KEYINPUT95), .B(n539), .Z(n376) );
  NOR2_X1 U449 ( .A1(n541), .A2(n376), .ZN(n377) );
  XNOR2_X1 U450 ( .A(n377), .B(KEYINPUT96), .ZN(n378) );
  NOR2_X1 U451 ( .A1(n379), .A2(n378), .ZN(n500) );
  XOR2_X1 U452 ( .A(KEYINPUT14), .B(KEYINPUT78), .Z(n381) );
  XNOR2_X1 U453 ( .A(KEYINPUT12), .B(KEYINPUT79), .ZN(n380) );
  XNOR2_X1 U454 ( .A(n381), .B(n380), .ZN(n386) );
  XOR2_X1 U455 ( .A(G57GAT), .B(KEYINPUT13), .Z(n427) );
  XOR2_X1 U456 ( .A(n427), .B(G71GAT), .Z(n384) );
  XNOR2_X1 U457 ( .A(G183GAT), .B(n382), .ZN(n383) );
  XNOR2_X1 U458 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U459 ( .A(n386), .B(n385), .Z(n388) );
  NAND2_X1 U460 ( .A1(G231GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U461 ( .A(n388), .B(n387), .ZN(n396) );
  XOR2_X1 U462 ( .A(G211GAT), .B(G78GAT), .Z(n390) );
  XNOR2_X1 U463 ( .A(G22GAT), .B(G155GAT), .ZN(n389) );
  XNOR2_X1 U464 ( .A(n390), .B(n389), .ZN(n394) );
  XOR2_X1 U465 ( .A(KEYINPUT15), .B(G64GAT), .Z(n392) );
  XNOR2_X1 U466 ( .A(G1GAT), .B(G8GAT), .ZN(n391) );
  XNOR2_X1 U467 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U468 ( .A(n394), .B(n393), .Z(n395) );
  XNOR2_X1 U469 ( .A(n396), .B(n395), .ZN(n562) );
  NOR2_X1 U470 ( .A1(n500), .A2(n562), .ZN(n397) );
  XNOR2_X1 U471 ( .A(KEYINPUT104), .B(n397), .ZN(n418) );
  XOR2_X1 U472 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n399) );
  XNOR2_X1 U473 ( .A(G43GAT), .B(G29GAT), .ZN(n398) );
  XNOR2_X1 U474 ( .A(n399), .B(n398), .ZN(n400) );
  XOR2_X1 U475 ( .A(KEYINPUT71), .B(n400), .Z(n451) );
  XOR2_X1 U476 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n402) );
  XNOR2_X1 U477 ( .A(KEYINPUT65), .B(KEYINPUT9), .ZN(n401) );
  XNOR2_X1 U478 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U479 ( .A(n451), .B(n403), .ZN(n417) );
  NAND2_X1 U480 ( .A1(G232GAT), .A2(G233GAT), .ZN(n405) );
  INV_X1 U481 ( .A(KEYINPUT11), .ZN(n404) );
  XOR2_X1 U482 ( .A(G92GAT), .B(G85GAT), .Z(n409) );
  XNOR2_X1 U483 ( .A(G99GAT), .B(G106GAT), .ZN(n408) );
  XNOR2_X1 U484 ( .A(n409), .B(n408), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U486 ( .A(n566), .B(KEYINPUT77), .ZN(n569) );
  XOR2_X1 U487 ( .A(KEYINPUT36), .B(n569), .Z(n589) );
  AND2_X1 U488 ( .A1(n418), .A2(n589), .ZN(n419) );
  XNOR2_X1 U489 ( .A(KEYINPUT37), .B(n419), .ZN(n485) );
  XOR2_X1 U490 ( .A(KEYINPUT75), .B(KEYINPUT72), .Z(n421) );
  XNOR2_X1 U491 ( .A(KEYINPUT73), .B(KEYINPUT33), .ZN(n420) );
  XNOR2_X1 U492 ( .A(n421), .B(n420), .ZN(n434) );
  NAND2_X1 U493 ( .A1(G230GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U494 ( .A(n295), .B(n424), .ZN(n425) );
  XOR2_X1 U495 ( .A(n425), .B(KEYINPUT32), .Z(n432) );
  XNOR2_X1 U496 ( .A(n426), .B(KEYINPUT31), .ZN(n430) );
  XNOR2_X1 U497 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n458) );
  INV_X1 U499 ( .A(n458), .ZN(n583) );
  XOR2_X1 U500 ( .A(KEYINPUT108), .B(n557), .Z(n543) );
  XOR2_X1 U501 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n436) );
  NAND2_X1 U502 ( .A1(G229GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U503 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U504 ( .A(KEYINPUT70), .B(n437), .ZN(n449) );
  XOR2_X1 U505 ( .A(G113GAT), .B(G15GAT), .Z(n441) );
  XNOR2_X1 U506 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U507 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U508 ( .A(n442), .B(G36GAT), .Z(n447) );
  XOR2_X1 U509 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n444) );
  XNOR2_X1 U510 ( .A(G197GAT), .B(G1GAT), .ZN(n443) );
  XNOR2_X1 U511 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U512 ( .A(n445), .B(G50GAT), .ZN(n446) );
  XNOR2_X1 U513 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U514 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U515 ( .A(n451), .B(n450), .ZN(n578) );
  INV_X1 U516 ( .A(n578), .ZN(n555) );
  OR2_X1 U517 ( .A1(n543), .A2(n555), .ZN(n520) );
  NOR2_X1 U518 ( .A1(n485), .A2(n520), .ZN(n535) );
  NAND2_X1 U519 ( .A1(n527), .A2(n535), .ZN(n453) );
  XNOR2_X1 U520 ( .A(n453), .B(n452), .ZN(G1339GAT) );
  NAND2_X1 U521 ( .A1(n523), .A2(n535), .ZN(n455) );
  INV_X1 U522 ( .A(KEYINPUT115), .ZN(n464) );
  NAND2_X1 U523 ( .A1(n562), .A2(n589), .ZN(n457) );
  XNOR2_X1 U524 ( .A(n457), .B(n456), .ZN(n459) );
  NOR2_X1 U525 ( .A1(n459), .A2(n458), .ZN(n461) );
  INV_X1 U526 ( .A(KEYINPUT114), .ZN(n460) );
  XNOR2_X1 U527 ( .A(n461), .B(n460), .ZN(n462) );
  NOR2_X1 U528 ( .A1(n462), .A2(n555), .ZN(n463) );
  XNOR2_X1 U529 ( .A(n464), .B(n463), .ZN(n470) );
  NAND2_X1 U530 ( .A1(n555), .A2(n557), .ZN(n465) );
  XNOR2_X1 U531 ( .A(KEYINPUT46), .B(n465), .ZN(n467) );
  INV_X1 U532 ( .A(n562), .ZN(n586) );
  NOR2_X1 U533 ( .A1(n562), .A2(n566), .ZN(n466) );
  XOR2_X1 U534 ( .A(KEYINPUT47), .B(n468), .Z(n469) );
  NOR2_X1 U535 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U536 ( .A(n471), .B(KEYINPUT48), .ZN(n538) );
  NOR2_X1 U537 ( .A1(n472), .A2(n538), .ZN(n474) );
  INV_X1 U538 ( .A(KEYINPUT54), .ZN(n473) );
  XNOR2_X1 U539 ( .A(n474), .B(n473), .ZN(n475) );
  NOR2_X1 U540 ( .A1(n475), .A2(n532), .ZN(n577) );
  NAND2_X1 U541 ( .A1(n577), .A2(n476), .ZN(n477) );
  XNOR2_X1 U542 ( .A(n477), .B(KEYINPUT55), .ZN(n478) );
  NAND2_X1 U543 ( .A1(n478), .A2(n541), .ZN(n482) );
  NOR2_X1 U544 ( .A1(n482), .A2(n543), .ZN(n481) );
  XNOR2_X1 U545 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n479) );
  XNOR2_X1 U546 ( .A(n479), .B(G176GAT), .ZN(n480) );
  XNOR2_X1 U547 ( .A(n481), .B(n480), .ZN(G1349GAT) );
  NOR2_X1 U548 ( .A1(n578), .A2(n482), .ZN(n484) );
  XNOR2_X1 U549 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n483) );
  XNOR2_X1 U550 ( .A(n484), .B(n483), .ZN(G1348GAT) );
  NAND2_X1 U551 ( .A1(n555), .A2(n583), .ZN(n503) );
  AND2_X1 U552 ( .A1(n532), .A2(n516), .ZN(n490) );
  XNOR2_X1 U553 ( .A(KEYINPUT105), .B(KEYINPUT39), .ZN(n488) );
  XNOR2_X1 U554 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U555 ( .A(n490), .B(n489), .ZN(G1328GAT) );
  AND2_X1 U556 ( .A1(n541), .A2(n516), .ZN(n494) );
  XNOR2_X1 U557 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n492) );
  XNOR2_X1 U558 ( .A(n494), .B(n493), .ZN(G1330GAT) );
  NOR2_X1 U559 ( .A1(n586), .A2(n482), .ZN(n497) );
  INV_X1 U560 ( .A(G183GAT), .ZN(n495) );
  XOR2_X1 U561 ( .A(KEYINPUT34), .B(KEYINPUT100), .Z(n505) );
  XOR2_X1 U562 ( .A(KEYINPUT16), .B(KEYINPUT80), .Z(n499) );
  NAND2_X1 U563 ( .A1(n569), .A2(n562), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(n502) );
  INV_X1 U565 ( .A(n500), .ZN(n501) );
  NAND2_X1 U566 ( .A1(n502), .A2(n501), .ZN(n519) );
  NOR2_X1 U567 ( .A1(n503), .A2(n519), .ZN(n512) );
  NAND2_X1 U568 ( .A1(n512), .A2(n532), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U570 ( .A(G1GAT), .B(n506), .Z(G1324GAT) );
  NAND2_X1 U571 ( .A1(n523), .A2(n512), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n507), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n509) );
  NAND2_X1 U574 ( .A1(n512), .A2(n541), .ZN(n508) );
  XNOR2_X1 U575 ( .A(n509), .B(n508), .ZN(n511) );
  XOR2_X1 U576 ( .A(G15GAT), .B(KEYINPUT101), .Z(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(G1326GAT) );
  XOR2_X1 U578 ( .A(G22GAT), .B(KEYINPUT103), .Z(n514) );
  NAND2_X1 U579 ( .A1(n512), .A2(n527), .ZN(n513) );
  XNOR2_X1 U580 ( .A(n514), .B(n513), .ZN(G1327GAT) );
  NAND2_X1 U581 ( .A1(n516), .A2(n523), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n515), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U583 ( .A(G50GAT), .B(KEYINPUT107), .Z(n518) );
  NAND2_X1 U584 ( .A1(n516), .A2(n527), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(G1331GAT) );
  XNOR2_X1 U586 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n522) );
  NOR2_X1 U587 ( .A1(n520), .A2(n519), .ZN(n528) );
  NAND2_X1 U588 ( .A1(n532), .A2(n528), .ZN(n521) );
  XNOR2_X1 U589 ( .A(n522), .B(n521), .ZN(G1332GAT) );
  NAND2_X1 U590 ( .A1(n523), .A2(n528), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U592 ( .A(G71GAT), .B(KEYINPUT109), .Z(n526) );
  NAND2_X1 U593 ( .A1(n528), .A2(n541), .ZN(n525) );
  XNOR2_X1 U594 ( .A(n526), .B(n525), .ZN(G1334GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n530) );
  NAND2_X1 U596 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(G78GAT), .B(n531), .ZN(G1335GAT) );
  XOR2_X1 U599 ( .A(G85GAT), .B(KEYINPUT111), .Z(n534) );
  NAND2_X1 U600 ( .A1(n535), .A2(n532), .ZN(n533) );
  XNOR2_X1 U601 ( .A(n534), .B(n533), .ZN(G1336GAT) );
  XOR2_X1 U602 ( .A(G99GAT), .B(KEYINPUT113), .Z(n537) );
  NAND2_X1 U603 ( .A1(n535), .A2(n541), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(G1338GAT) );
  NOR2_X1 U605 ( .A1(n538), .A2(n539), .ZN(n540) );
  NAND2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n549) );
  NOR2_X1 U607 ( .A1(n578), .A2(n549), .ZN(n542) );
  XOR2_X1 U608 ( .A(G113GAT), .B(n542), .Z(G1340GAT) );
  NOR2_X1 U609 ( .A1(n543), .A2(n549), .ZN(n545) );
  XNOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(G1341GAT) );
  NOR2_X1 U612 ( .A1(n586), .A2(n549), .ZN(n547) );
  XNOR2_X1 U613 ( .A(KEYINPUT116), .B(KEYINPUT50), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U615 ( .A(G127GAT), .B(n548), .Z(G1342GAT) );
  NOR2_X1 U616 ( .A1(n569), .A2(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(n552) );
  XOR2_X1 U619 ( .A(G134GAT), .B(n552), .Z(G1343GAT) );
  NAND2_X1 U620 ( .A1(n576), .A2(n553), .ZN(n554) );
  NOR2_X1 U621 ( .A1(n538), .A2(n554), .ZN(n565) );
  NAND2_X1 U622 ( .A1(n565), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n561) );
  XOR2_X1 U625 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n559) );
  NAND2_X1 U626 ( .A1(n565), .A2(n557), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1345GAT) );
  XOR2_X1 U629 ( .A(G155GAT), .B(KEYINPUT119), .Z(n564) );
  NAND2_X1 U630 ( .A1(n565), .A2(n562), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1346GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(KEYINPUT120), .ZN(n568) );
  XNOR2_X1 U634 ( .A(G162GAT), .B(n568), .ZN(G1347GAT) );
  NOR2_X1 U635 ( .A1(n482), .A2(n569), .ZN(n573) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(KEYINPUT123), .ZN(n571) );
  XNOR2_X1 U638 ( .A(KEYINPUT124), .B(n571), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(G1351GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT127), .B(KEYINPUT126), .Z(n575) );
  XNOR2_X1 U641 ( .A(KEYINPUT125), .B(KEYINPUT60), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(n582) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n588) );
  NOR2_X1 U644 ( .A1(n578), .A2(n588), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n581) );
  XOR2_X1 U647 ( .A(n582), .B(n581), .Z(G1352GAT) );
  NOR2_X1 U648 ( .A1(n583), .A2(n588), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1353GAT) );
  NOR2_X1 U651 ( .A1(n586), .A2(n588), .ZN(n587) );
  XOR2_X1 U652 ( .A(G211GAT), .B(n587), .Z(G1354GAT) );
  INV_X1 U653 ( .A(n588), .ZN(n590) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(KEYINPUT62), .ZN(n592) );
  XNOR2_X1 U656 ( .A(G218GAT), .B(n592), .ZN(G1355GAT) );
endmodule

