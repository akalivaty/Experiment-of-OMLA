

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598;

  NOR2_X1 U323 ( .A1(n472), .A2(n471), .ZN(n475) );
  XOR2_X1 U324 ( .A(G36GAT), .B(G218GAT), .Z(n430) );
  XNOR2_X1 U325 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U326 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U327 ( .A(n439), .B(n438), .ZN(n443) );
  XNOR2_X1 U328 ( .A(n437), .B(n293), .ZN(n438) );
  XNOR2_X1 U329 ( .A(n365), .B(n364), .ZN(n369) );
  XNOR2_X1 U330 ( .A(n451), .B(n450), .ZN(n532) );
  XNOR2_X1 U331 ( .A(n449), .B(KEYINPUT102), .ZN(n450) );
  INV_X1 U332 ( .A(KEYINPUT37), .ZN(n449) );
  XOR2_X1 U333 ( .A(n370), .B(n415), .Z(n291) );
  AND2_X1 U334 ( .A1(G226GAT), .A2(G233GAT), .ZN(n292) );
  XOR2_X1 U335 ( .A(n436), .B(n435), .Z(n293) );
  XNOR2_X1 U336 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n459) );
  XNOR2_X1 U337 ( .A(KEYINPUT114), .B(KEYINPUT45), .ZN(n466) );
  XNOR2_X1 U338 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U339 ( .A(n414), .B(n312), .ZN(n313) );
  XNOR2_X1 U340 ( .A(n314), .B(n313), .ZN(n316) );
  INV_X1 U341 ( .A(KEYINPUT48), .ZN(n473) );
  XNOR2_X1 U342 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n476) );
  XNOR2_X1 U343 ( .A(n473), .B(KEYINPUT64), .ZN(n474) );
  XNOR2_X1 U344 ( .A(n323), .B(n336), .ZN(n324) );
  XNOR2_X1 U345 ( .A(n475), .B(n474), .ZN(n545) );
  XNOR2_X1 U346 ( .A(n430), .B(n292), .ZN(n364) );
  XNOR2_X1 U347 ( .A(n325), .B(n324), .ZN(n327) );
  NOR2_X1 U348 ( .A1(n533), .A2(n478), .ZN(n578) );
  XNOR2_X1 U349 ( .A(n371), .B(n291), .ZN(n372) );
  XNOR2_X1 U350 ( .A(KEYINPUT38), .B(KEYINPUT103), .ZN(n452) );
  XNOR2_X1 U351 ( .A(n447), .B(n446), .ZN(n574) );
  XNOR2_X1 U352 ( .A(n373), .B(n372), .ZN(n535) );
  XNOR2_X1 U353 ( .A(n453), .B(n452), .ZN(n515) );
  XNOR2_X1 U354 ( .A(n487), .B(G176GAT), .ZN(n488) );
  XNOR2_X1 U355 ( .A(n455), .B(G36GAT), .ZN(n456) );
  XNOR2_X1 U356 ( .A(n489), .B(n488), .ZN(G1349GAT) );
  XNOR2_X1 U357 ( .A(n457), .B(n456), .ZN(G1329GAT) );
  XOR2_X1 U358 ( .A(G1GAT), .B(G141GAT), .Z(n295) );
  XNOR2_X1 U359 ( .A(G169GAT), .B(G197GAT), .ZN(n294) );
  XNOR2_X1 U360 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U361 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n297) );
  XNOR2_X1 U362 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n296) );
  XNOR2_X1 U363 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U364 ( .A(n299), .B(n298), .ZN(n310) );
  XNOR2_X1 U365 ( .A(G113GAT), .B(G15GAT), .ZN(n360) );
  XOR2_X1 U366 ( .A(G22GAT), .B(G50GAT), .Z(n301) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(G36GAT), .ZN(n300) );
  XNOR2_X1 U368 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U369 ( .A(n360), .B(n302), .ZN(n304) );
  NAND2_X1 U370 ( .A1(G229GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U371 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U372 ( .A(n305), .B(KEYINPUT67), .Z(n308) );
  XNOR2_X1 U373 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n306) );
  XNOR2_X1 U374 ( .A(n306), .B(KEYINPUT7), .ZN(n445) );
  XNOR2_X1 U375 ( .A(n445), .B(KEYINPUT68), .ZN(n307) );
  XNOR2_X1 U376 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U377 ( .A(n310), .B(n309), .Z(n517) );
  INV_X1 U378 ( .A(n517), .ZN(n581) );
  XNOR2_X1 U379 ( .A(KEYINPUT70), .B(KEYINPUT32), .ZN(n311) );
  XOR2_X1 U380 ( .A(G176GAT), .B(G64GAT), .Z(n370) );
  XNOR2_X1 U381 ( .A(n311), .B(n370), .ZN(n314) );
  XOR2_X1 U382 ( .A(G57GAT), .B(KEYINPUT13), .Z(n414) );
  AND2_X1 U383 ( .A1(G230GAT), .A2(G233GAT), .ZN(n312) );
  INV_X1 U384 ( .A(KEYINPUT33), .ZN(n315) );
  NAND2_X1 U385 ( .A1(n316), .A2(n315), .ZN(n319) );
  INV_X1 U386 ( .A(n316), .ZN(n317) );
  NAND2_X1 U387 ( .A1(n317), .A2(KEYINPUT33), .ZN(n318) );
  NAND2_X1 U388 ( .A1(n319), .A2(n318), .ZN(n325) );
  XNOR2_X1 U389 ( .A(G85GAT), .B(KEYINPUT69), .ZN(n320) );
  XNOR2_X1 U390 ( .A(n320), .B(G92GAT), .ZN(n444) );
  XNOR2_X1 U391 ( .A(n444), .B(KEYINPUT31), .ZN(n323) );
  XOR2_X1 U392 ( .A(G78GAT), .B(G148GAT), .Z(n322) );
  XNOR2_X1 U393 ( .A(G106GAT), .B(G204GAT), .ZN(n321) );
  XNOR2_X1 U394 ( .A(n322), .B(n321), .ZN(n336) );
  XOR2_X1 U395 ( .A(G99GAT), .B(G71GAT), .Z(n326) );
  XOR2_X1 U396 ( .A(G120GAT), .B(n326), .Z(n353) );
  XNOR2_X1 U397 ( .A(n327), .B(n353), .ZN(n586) );
  INV_X1 U398 ( .A(n586), .ZN(n328) );
  NAND2_X1 U399 ( .A1(n581), .A2(n328), .ZN(n495) );
  XOR2_X1 U400 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n330) );
  XNOR2_X1 U401 ( .A(G218GAT), .B(KEYINPUT81), .ZN(n329) );
  XNOR2_X1 U402 ( .A(n330), .B(n329), .ZN(n345) );
  XOR2_X1 U403 ( .A(KEYINPUT84), .B(KEYINPUT24), .Z(n332) );
  NAND2_X1 U404 ( .A1(G228GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U405 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U406 ( .A(n333), .B(KEYINPUT85), .Z(n338) );
  XOR2_X1 U407 ( .A(G211GAT), .B(KEYINPUT82), .Z(n335) );
  XNOR2_X1 U408 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n334) );
  XNOR2_X1 U409 ( .A(n335), .B(n334), .ZN(n365) );
  XNOR2_X1 U410 ( .A(n365), .B(n336), .ZN(n337) );
  XNOR2_X1 U411 ( .A(n338), .B(n337), .ZN(n341) );
  XOR2_X1 U412 ( .A(KEYINPUT83), .B(KEYINPUT3), .Z(n340) );
  XNOR2_X1 U413 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n339) );
  XNOR2_X1 U414 ( .A(n340), .B(n339), .ZN(n383) );
  XOR2_X1 U415 ( .A(n341), .B(n383), .Z(n343) );
  XOR2_X1 U416 ( .A(G50GAT), .B(G162GAT), .Z(n431) );
  XOR2_X1 U417 ( .A(G22GAT), .B(G155GAT), .Z(n425) );
  XNOR2_X1 U418 ( .A(n431), .B(n425), .ZN(n342) );
  XNOR2_X1 U419 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U420 ( .A(n345), .B(n344), .Z(n479) );
  XNOR2_X1 U421 ( .A(n479), .B(KEYINPUT28), .ZN(n514) );
  INV_X1 U422 ( .A(n514), .ZN(n550) );
  XNOR2_X1 U423 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n346) );
  XNOR2_X1 U424 ( .A(n346), .B(KEYINPUT19), .ZN(n347) );
  XOR2_X1 U425 ( .A(n347), .B(KEYINPUT17), .Z(n349) );
  XNOR2_X1 U426 ( .A(G169GAT), .B(G190GAT), .ZN(n348) );
  XNOR2_X1 U427 ( .A(n349), .B(n348), .ZN(n371) );
  XOR2_X1 U428 ( .A(KEYINPUT78), .B(KEYINPUT20), .Z(n351) );
  XNOR2_X1 U429 ( .A(KEYINPUT79), .B(KEYINPUT76), .ZN(n350) );
  XNOR2_X1 U430 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U431 ( .A(n371), .B(n352), .ZN(n363) );
  XOR2_X1 U432 ( .A(n353), .B(KEYINPUT77), .Z(n355) );
  NAND2_X1 U433 ( .A1(G227GAT), .A2(G233GAT), .ZN(n354) );
  XNOR2_X1 U434 ( .A(n355), .B(n354), .ZN(n359) );
  XOR2_X1 U435 ( .A(KEYINPUT75), .B(G176GAT), .Z(n357) );
  XOR2_X1 U436 ( .A(G43GAT), .B(G134GAT), .Z(n434) );
  XOR2_X1 U437 ( .A(KEYINPUT0), .B(G127GAT), .Z(n379) );
  XNOR2_X1 U438 ( .A(n434), .B(n379), .ZN(n356) );
  XNOR2_X1 U439 ( .A(n357), .B(n356), .ZN(n358) );
  XNOR2_X1 U440 ( .A(n359), .B(n358), .ZN(n361) );
  XNOR2_X1 U441 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U442 ( .A(n363), .B(n362), .Z(n547) );
  INV_X1 U443 ( .A(n547), .ZN(n539) );
  XOR2_X1 U444 ( .A(n539), .B(KEYINPUT80), .Z(n398) );
  INV_X1 U445 ( .A(G92GAT), .ZN(n374) );
  XOR2_X1 U446 ( .A(KEYINPUT90), .B(KEYINPUT92), .Z(n367) );
  XNOR2_X1 U447 ( .A(G204GAT), .B(KEYINPUT91), .ZN(n366) );
  XNOR2_X1 U448 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U449 ( .A(n369), .B(n368), .Z(n373) );
  XOR2_X1 U450 ( .A(G8GAT), .B(KEYINPUT73), .Z(n415) );
  XNOR2_X1 U451 ( .A(n374), .B(n535), .ZN(n522) );
  INV_X1 U452 ( .A(n522), .ZN(n454) );
  XOR2_X1 U453 ( .A(n454), .B(KEYINPUT93), .Z(n375) );
  XNOR2_X1 U454 ( .A(n375), .B(KEYINPUT27), .ZN(n402) );
  XOR2_X1 U455 ( .A(G85GAT), .B(G162GAT), .Z(n377) );
  XNOR2_X1 U456 ( .A(G29GAT), .B(G134GAT), .ZN(n376) );
  XNOR2_X1 U457 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U458 ( .A(n379), .B(n378), .Z(n381) );
  NAND2_X1 U459 ( .A1(G225GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U460 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U461 ( .A(n382), .B(KEYINPUT86), .Z(n385) );
  XNOR2_X1 U462 ( .A(n383), .B(KEYINPUT88), .ZN(n384) );
  XNOR2_X1 U463 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U464 ( .A(G155GAT), .B(G148GAT), .Z(n387) );
  XNOR2_X1 U465 ( .A(G113GAT), .B(G120GAT), .ZN(n386) );
  XNOR2_X1 U466 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U467 ( .A(n389), .B(n388), .Z(n397) );
  XOR2_X1 U468 ( .A(KEYINPUT1), .B(KEYINPUT89), .Z(n391) );
  XNOR2_X1 U469 ( .A(G57GAT), .B(KEYINPUT6), .ZN(n390) );
  XNOR2_X1 U470 ( .A(n391), .B(n390), .ZN(n395) );
  XOR2_X1 U471 ( .A(KEYINPUT87), .B(KEYINPUT4), .Z(n393) );
  XNOR2_X1 U472 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n392) );
  XNOR2_X1 U473 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U474 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U475 ( .A(n397), .B(n396), .Z(n508) );
  NOR2_X1 U476 ( .A1(n402), .A2(n508), .ZN(n546) );
  NAND2_X1 U477 ( .A1(n398), .A2(n546), .ZN(n399) );
  NOR2_X1 U478 ( .A1(n550), .A2(n399), .ZN(n400) );
  XNOR2_X1 U479 ( .A(n400), .B(KEYINPUT94), .ZN(n411) );
  INV_X1 U480 ( .A(n508), .ZN(n533) );
  NOR2_X1 U481 ( .A1(n539), .A2(n479), .ZN(n401) );
  XOR2_X1 U482 ( .A(n401), .B(KEYINPUT26), .Z(n579) );
  NOR2_X1 U483 ( .A1(n402), .A2(n579), .ZN(n403) );
  XOR2_X1 U484 ( .A(KEYINPUT95), .B(n403), .Z(n408) );
  NAND2_X1 U485 ( .A1(n539), .A2(n522), .ZN(n404) );
  NAND2_X1 U486 ( .A1(n404), .A2(n479), .ZN(n405) );
  XNOR2_X1 U487 ( .A(n405), .B(KEYINPUT96), .ZN(n406) );
  XNOR2_X1 U488 ( .A(KEYINPUT25), .B(n406), .ZN(n407) );
  NOR2_X1 U489 ( .A1(n408), .A2(n407), .ZN(n409) );
  NOR2_X1 U490 ( .A1(n533), .A2(n409), .ZN(n410) );
  NOR2_X1 U491 ( .A1(n411), .A2(n410), .ZN(n492) );
  XOR2_X1 U492 ( .A(G78GAT), .B(G211GAT), .Z(n413) );
  XNOR2_X1 U493 ( .A(G15GAT), .B(G127GAT), .ZN(n412) );
  XNOR2_X1 U494 ( .A(n413), .B(n412), .ZN(n429) );
  XOR2_X1 U495 ( .A(n415), .B(n414), .Z(n417) );
  NAND2_X1 U496 ( .A1(G231GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U497 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U498 ( .A(KEYINPUT15), .B(KEYINPUT74), .Z(n419) );
  XNOR2_X1 U499 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n418) );
  XNOR2_X1 U500 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U501 ( .A(n421), .B(n420), .Z(n427) );
  XOR2_X1 U502 ( .A(G64GAT), .B(G71GAT), .Z(n423) );
  XNOR2_X1 U503 ( .A(G1GAT), .B(G183GAT), .ZN(n422) );
  XNOR2_X1 U504 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U505 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U506 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U507 ( .A(n429), .B(n428), .ZN(n591) );
  NOR2_X1 U508 ( .A1(n492), .A2(n591), .ZN(n448) );
  XOR2_X1 U509 ( .A(KEYINPUT9), .B(KEYINPUT65), .Z(n433) );
  XNOR2_X1 U510 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U511 ( .A(n433), .B(n432), .ZN(n439) );
  XNOR2_X1 U512 ( .A(G190GAT), .B(n434), .ZN(n437) );
  XOR2_X1 U513 ( .A(KEYINPUT10), .B(G99GAT), .Z(n436) );
  NAND2_X1 U514 ( .A1(G232GAT), .A2(G233GAT), .ZN(n435) );
  XOR2_X1 U515 ( .A(KEYINPUT72), .B(KEYINPUT11), .Z(n441) );
  XNOR2_X1 U516 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n440) );
  XNOR2_X1 U517 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U518 ( .A(n443), .B(n442), .ZN(n447) );
  XNOR2_X1 U519 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U520 ( .A(KEYINPUT36), .B(n574), .ZN(n594) );
  NAND2_X1 U521 ( .A1(n448), .A2(n594), .ZN(n451) );
  NOR2_X1 U522 ( .A1(n495), .A2(n532), .ZN(n453) );
  NOR2_X1 U523 ( .A1(n515), .A2(n454), .ZN(n457) );
  INV_X1 U524 ( .A(KEYINPUT104), .ZN(n455) );
  INV_X1 U525 ( .A(KEYINPUT41), .ZN(n458) );
  XNOR2_X1 U526 ( .A(n458), .B(n586), .ZN(n564) );
  NAND2_X1 U527 ( .A1(n564), .A2(n581), .ZN(n460) );
  INV_X1 U528 ( .A(n591), .ZN(n490) );
  NAND2_X1 U529 ( .A1(n461), .A2(n490), .ZN(n462) );
  XNOR2_X1 U530 ( .A(n462), .B(KEYINPUT113), .ZN(n464) );
  INV_X1 U531 ( .A(n574), .ZN(n463) );
  NAND2_X1 U532 ( .A1(n464), .A2(n463), .ZN(n465) );
  XNOR2_X1 U533 ( .A(n465), .B(KEYINPUT47), .ZN(n472) );
  NAND2_X1 U534 ( .A1(n594), .A2(n591), .ZN(n467) );
  NOR2_X1 U535 ( .A1(n468), .A2(n586), .ZN(n469) );
  XNOR2_X1 U536 ( .A(n469), .B(KEYINPUT115), .ZN(n470) );
  NOR2_X1 U537 ( .A1(n470), .A2(n581), .ZN(n471) );
  NAND2_X1 U538 ( .A1(n545), .A2(n522), .ZN(n477) );
  NAND2_X1 U539 ( .A1(n479), .A2(n578), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n480), .B(KEYINPUT55), .ZN(n481) );
  NAND2_X1 U541 ( .A1(n481), .A2(n539), .ZN(n484) );
  INV_X1 U542 ( .A(n484), .ZN(n483) );
  INV_X1 U543 ( .A(KEYINPUT121), .ZN(n482) );
  NAND2_X1 U544 ( .A1(n483), .A2(n482), .ZN(n486) );
  NAND2_X1 U545 ( .A1(KEYINPUT121), .A2(n484), .ZN(n485) );
  NAND2_X1 U546 ( .A1(n486), .A2(n485), .ZN(n575) );
  XNOR2_X1 U547 ( .A(n564), .B(KEYINPUT106), .ZN(n553) );
  NAND2_X1 U548 ( .A1(n575), .A2(n553), .ZN(n489) );
  XOR2_X1 U549 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n487) );
  NOR2_X1 U550 ( .A1(n490), .A2(n574), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n491), .B(KEYINPUT16), .ZN(n494) );
  INV_X1 U552 ( .A(n492), .ZN(n493) );
  NAND2_X1 U553 ( .A1(n494), .A2(n493), .ZN(n519) );
  NOR2_X1 U554 ( .A1(n495), .A2(n519), .ZN(n504) );
  NAND2_X1 U555 ( .A1(n504), .A2(n533), .ZN(n498) );
  XOR2_X1 U556 ( .A(G1GAT), .B(KEYINPUT97), .Z(n496) );
  XNOR2_X1 U557 ( .A(KEYINPUT34), .B(n496), .ZN(n497) );
  XNOR2_X1 U558 ( .A(n498), .B(n497), .ZN(G1324GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n500) );
  NAND2_X1 U560 ( .A1(n504), .A2(n522), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G8GAT), .B(n501), .ZN(G1325GAT) );
  XOR2_X1 U563 ( .A(G15GAT), .B(KEYINPUT35), .Z(n503) );
  NAND2_X1 U564 ( .A1(n504), .A2(n539), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(G1326GAT) );
  XOR2_X1 U566 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n506) );
  NAND2_X1 U567 ( .A1(n504), .A2(n550), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U569 ( .A(G22GAT), .B(n507), .ZN(G1327GAT) );
  NOR2_X1 U570 ( .A1(n515), .A2(n508), .ZN(n510) );
  XNOR2_X1 U571 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(G1328GAT) );
  XNOR2_X1 U573 ( .A(KEYINPUT105), .B(KEYINPUT40), .ZN(n512) );
  NOR2_X1 U574 ( .A1(n547), .A2(n515), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U576 ( .A(G43GAT), .B(n513), .ZN(G1330GAT) );
  NOR2_X1 U577 ( .A1(n515), .A2(n514), .ZN(n516) );
  XOR2_X1 U578 ( .A(G50GAT), .B(n516), .Z(G1331GAT) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n521) );
  NAND2_X1 U580 ( .A1(n553), .A2(n517), .ZN(n518) );
  XOR2_X1 U581 ( .A(KEYINPUT107), .B(n518), .Z(n531) );
  NOR2_X1 U582 ( .A1(n531), .A2(n519), .ZN(n528) );
  NAND2_X1 U583 ( .A1(n533), .A2(n528), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n521), .B(n520), .ZN(G1332GAT) );
  NAND2_X1 U585 ( .A1(n528), .A2(n522), .ZN(n523) );
  XNOR2_X1 U586 ( .A(n523), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U587 ( .A1(n539), .A2(n528), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n524), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n526) );
  XNOR2_X1 U590 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U592 ( .A(KEYINPUT108), .B(n527), .Z(n530) );
  NAND2_X1 U593 ( .A1(n528), .A2(n550), .ZN(n529) );
  XNOR2_X1 U594 ( .A(n530), .B(n529), .ZN(G1335GAT) );
  NOR2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n541) );
  NAND2_X1 U596 ( .A1(n541), .A2(n533), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n534), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U598 ( .A1(n535), .A2(n541), .ZN(n538) );
  INV_X1 U599 ( .A(n541), .ZN(n536) );
  NAND2_X1 U600 ( .A1(G92GAT), .A2(n536), .ZN(n537) );
  NAND2_X1 U601 ( .A1(n538), .A2(n537), .ZN(G1337GAT) );
  NAND2_X1 U602 ( .A1(n539), .A2(n541), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n540), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT111), .B(KEYINPUT44), .Z(n543) );
  NAND2_X1 U605 ( .A1(n541), .A2(n550), .ZN(n542) );
  XNOR2_X1 U606 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U607 ( .A(G106GAT), .B(n544), .ZN(G1339GAT) );
  XOR2_X1 U608 ( .A(G113GAT), .B(KEYINPUT117), .Z(n552) );
  NAND2_X1 U609 ( .A1(n546), .A2(n545), .ZN(n561) );
  NOR2_X1 U610 ( .A1(n547), .A2(n561), .ZN(n548) );
  XOR2_X1 U611 ( .A(KEYINPUT116), .B(n548), .Z(n549) );
  NOR2_X1 U612 ( .A1(n550), .A2(n549), .ZN(n558) );
  NAND2_X1 U613 ( .A1(n558), .A2(n581), .ZN(n551) );
  XNOR2_X1 U614 ( .A(n552), .B(n551), .ZN(G1340GAT) );
  XOR2_X1 U615 ( .A(G120GAT), .B(KEYINPUT49), .Z(n555) );
  NAND2_X1 U616 ( .A1(n558), .A2(n553), .ZN(n554) );
  XNOR2_X1 U617 ( .A(n555), .B(n554), .ZN(G1341GAT) );
  NAND2_X1 U618 ( .A1(n591), .A2(n558), .ZN(n556) );
  XNOR2_X1 U619 ( .A(n556), .B(KEYINPUT50), .ZN(n557) );
  XNOR2_X1 U620 ( .A(G127GAT), .B(n557), .ZN(G1342GAT) );
  XOR2_X1 U621 ( .A(G134GAT), .B(KEYINPUT51), .Z(n560) );
  NAND2_X1 U622 ( .A1(n558), .A2(n574), .ZN(n559) );
  XNOR2_X1 U623 ( .A(n560), .B(n559), .ZN(G1343GAT) );
  NOR2_X1 U624 ( .A1(n561), .A2(n579), .ZN(n562) );
  XNOR2_X1 U625 ( .A(n562), .B(KEYINPUT118), .ZN(n570) );
  NAND2_X1 U626 ( .A1(n570), .A2(n581), .ZN(n563) );
  XNOR2_X1 U627 ( .A(n563), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n566) );
  NAND2_X1 U629 ( .A1(n564), .A2(n570), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n566), .B(n565), .ZN(n568) );
  XOR2_X1 U631 ( .A(G148GAT), .B(KEYINPUT119), .Z(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(G1345GAT) );
  NAND2_X1 U633 ( .A1(n570), .A2(n591), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U635 ( .A1(n570), .A2(n574), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U637 ( .A1(n575), .A2(n581), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U639 ( .A1(n591), .A2(n575), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n573), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U641 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1351GAT) );
  INV_X1 U644 ( .A(n578), .ZN(n580) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n595) );
  NAND2_X1 U646 ( .A1(n595), .A2(n581), .ZN(n585) );
  XOR2_X1 U647 ( .A(KEYINPUT60), .B(KEYINPUT122), .Z(n583) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n582) );
  XNOR2_X1 U649 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT61), .B(KEYINPUT124), .Z(n588) );
  NAND2_X1 U652 ( .A1(n595), .A2(n586), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(n590) );
  XOR2_X1 U654 ( .A(G204GAT), .B(KEYINPUT123), .Z(n589) );
  XNOR2_X1 U655 ( .A(n590), .B(n589), .ZN(G1353GAT) );
  XOR2_X1 U656 ( .A(G211GAT), .B(KEYINPUT125), .Z(n593) );
  NAND2_X1 U657 ( .A1(n595), .A2(n591), .ZN(n592) );
  XNOR2_X1 U658 ( .A(n593), .B(n592), .ZN(G1354GAT) );
  XOR2_X1 U659 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n597) );
  NAND2_X1 U660 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U661 ( .A(n597), .B(n596), .ZN(n598) );
  XOR2_X1 U662 ( .A(G218GAT), .B(n598), .Z(G1355GAT) );
endmodule

