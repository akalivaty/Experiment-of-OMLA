

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580;

  XNOR2_X1 U321 ( .A(n361), .B(n306), .ZN(n307) );
  XNOR2_X1 U322 ( .A(n305), .B(n304), .ZN(n306) );
  INV_X1 U323 ( .A(G36GAT), .ZN(n304) );
  INV_X1 U324 ( .A(n517), .ZN(n472) );
  XNOR2_X1 U325 ( .A(n392), .B(n391), .ZN(n477) );
  XNOR2_X1 U326 ( .A(KEYINPUT97), .B(KEYINPUT96), .ZN(n366) );
  XOR2_X1 U327 ( .A(n474), .B(KEYINPUT28), .Z(n534) );
  INV_X1 U328 ( .A(n477), .ZN(n532) );
  XOR2_X1 U329 ( .A(n372), .B(n371), .Z(n289) );
  XOR2_X1 U330 ( .A(n461), .B(KEYINPUT47), .Z(n290) );
  XOR2_X1 U331 ( .A(n328), .B(n327), .Z(n291) );
  XOR2_X1 U332 ( .A(G120GAT), .B(KEYINPUT0), .Z(n292) );
  XOR2_X1 U333 ( .A(n428), .B(G15GAT), .Z(n293) );
  AND2_X1 U334 ( .A1(n473), .A2(n472), .ZN(n294) );
  XOR2_X1 U335 ( .A(n456), .B(KEYINPUT41), .Z(n546) );
  XNOR2_X1 U336 ( .A(KEYINPUT27), .B(KEYINPUT98), .ZN(n379) );
  XNOR2_X1 U337 ( .A(n520), .B(n379), .ZN(n443) );
  XNOR2_X1 U338 ( .A(n404), .B(n366), .ZN(n367) );
  INV_X1 U339 ( .A(G183GAT), .ZN(n385) );
  XNOR2_X1 U340 ( .A(KEYINPUT48), .B(KEYINPUT118), .ZN(n468) );
  XNOR2_X1 U341 ( .A(n386), .B(n385), .ZN(n387) );
  INV_X1 U342 ( .A(KEYINPUT66), .ZN(n311) );
  XNOR2_X1 U343 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U344 ( .A(n329), .B(n291), .ZN(n330) );
  XNOR2_X1 U345 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U346 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U347 ( .A(n314), .B(n313), .ZN(n315) );
  OR2_X1 U348 ( .A1(n490), .A2(n515), .ZN(n453) );
  XOR2_X1 U349 ( .A(KEYINPUT38), .B(n453), .Z(n503) );
  XNOR2_X1 U350 ( .A(n481), .B(G176GAT), .ZN(n482) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n454) );
  XNOR2_X1 U352 ( .A(n455), .B(n454), .ZN(G1330GAT) );
  XOR2_X1 U353 ( .A(KEYINPUT29), .B(KEYINPUT71), .Z(n296) );
  XNOR2_X1 U354 ( .A(KEYINPUT69), .B(KEYINPUT67), .ZN(n295) );
  XNOR2_X1 U355 ( .A(n296), .B(n295), .ZN(n316) );
  XOR2_X1 U356 ( .A(G197GAT), .B(G141GAT), .Z(n298) );
  XNOR2_X1 U357 ( .A(G169GAT), .B(G50GAT), .ZN(n297) );
  XNOR2_X1 U358 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U359 ( .A(KEYINPUT68), .B(G8GAT), .Z(n300) );
  XNOR2_X1 U360 ( .A(G113GAT), .B(G1GAT), .ZN(n299) );
  XNOR2_X1 U361 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U362 ( .A(n302), .B(n301), .Z(n309) );
  XNOR2_X1 U363 ( .A(G22GAT), .B(G15GAT), .ZN(n303) );
  XNOR2_X1 U364 ( .A(n303), .B(KEYINPUT70), .ZN(n361) );
  NAND2_X1 U365 ( .A1(G229GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U366 ( .A(G43GAT), .B(n307), .ZN(n308) );
  XNOR2_X1 U367 ( .A(n309), .B(n308), .ZN(n314) );
  XNOR2_X1 U368 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n310) );
  XNOR2_X1 U369 ( .A(n310), .B(KEYINPUT8), .ZN(n337) );
  XNOR2_X1 U370 ( .A(n337), .B(KEYINPUT30), .ZN(n312) );
  XOR2_X1 U371 ( .A(n316), .B(n315), .Z(n566) );
  INV_X1 U372 ( .A(n566), .ZN(n555) );
  XOR2_X1 U373 ( .A(G78GAT), .B(G148GAT), .Z(n318) );
  XNOR2_X1 U374 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n318), .B(n317), .ZN(n406) );
  XNOR2_X1 U376 ( .A(G71GAT), .B(G57GAT), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n319), .B(KEYINPUT13), .ZN(n355) );
  XOR2_X1 U378 ( .A(n406), .B(n355), .Z(n333) );
  XOR2_X1 U379 ( .A(G64GAT), .B(KEYINPUT76), .Z(n321) );
  XNOR2_X1 U380 ( .A(G204GAT), .B(G92GAT), .ZN(n320) );
  XNOR2_X1 U381 ( .A(n321), .B(n320), .ZN(n377) );
  XOR2_X1 U382 ( .A(G99GAT), .B(G85GAT), .Z(n334) );
  XOR2_X1 U383 ( .A(n377), .B(n334), .Z(n323) );
  XNOR2_X1 U384 ( .A(G176GAT), .B(G120GAT), .ZN(n322) );
  XNOR2_X1 U385 ( .A(n323), .B(n322), .ZN(n331) );
  XOR2_X1 U386 ( .A(KEYINPUT73), .B(KEYINPUT77), .Z(n325) );
  XNOR2_X1 U387 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n324) );
  XNOR2_X1 U388 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n326), .B(KEYINPUT72), .ZN(n329) );
  XOR2_X1 U390 ( .A(KEYINPUT32), .B(KEYINPUT75), .Z(n328) );
  NAND2_X1 U391 ( .A1(G230GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n569) );
  NAND2_X1 U393 ( .A1(n555), .A2(n569), .ZN(n490) );
  XOR2_X1 U394 ( .A(G36GAT), .B(G218GAT), .Z(n368) );
  XOR2_X1 U395 ( .A(n368), .B(n334), .Z(n336) );
  XOR2_X1 U396 ( .A(G43GAT), .B(G134GAT), .Z(n384) );
  XOR2_X1 U397 ( .A(G50GAT), .B(KEYINPUT78), .Z(n407) );
  XNOR2_X1 U398 ( .A(n384), .B(n407), .ZN(n335) );
  XNOR2_X1 U399 ( .A(n336), .B(n335), .ZN(n341) );
  XOR2_X1 U400 ( .A(G92GAT), .B(n337), .Z(n339) );
  NAND2_X1 U401 ( .A1(G232GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U402 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U403 ( .A(n341), .B(n340), .Z(n349) );
  XOR2_X1 U404 ( .A(KEYINPUT79), .B(KEYINPUT10), .Z(n343) );
  XNOR2_X1 U405 ( .A(KEYINPUT65), .B(KEYINPUT11), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U407 ( .A(KEYINPUT9), .B(G106GAT), .Z(n345) );
  XNOR2_X1 U408 ( .A(G190GAT), .B(G162GAT), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U410 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U411 ( .A(n349), .B(n348), .Z(n559) );
  XOR2_X1 U412 ( .A(KEYINPUT36), .B(n559), .Z(n578) );
  XOR2_X1 U413 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n351) );
  XNOR2_X1 U414 ( .A(G64GAT), .B(KEYINPUT80), .ZN(n350) );
  XOR2_X1 U415 ( .A(n351), .B(n350), .Z(n365) );
  XNOR2_X1 U416 ( .A(G8GAT), .B(G183GAT), .ZN(n352) );
  XNOR2_X1 U417 ( .A(n352), .B(G211GAT), .ZN(n371) );
  XOR2_X1 U418 ( .A(KEYINPUT81), .B(n371), .Z(n354) );
  NAND2_X1 U419 ( .A1(G231GAT), .A2(G233GAT), .ZN(n353) );
  XNOR2_X1 U420 ( .A(n354), .B(n353), .ZN(n356) );
  XOR2_X1 U421 ( .A(n356), .B(n355), .Z(n359) );
  XNOR2_X1 U422 ( .A(G1GAT), .B(G127GAT), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n357), .B(G155GAT), .ZN(n427) );
  XNOR2_X1 U424 ( .A(G78GAT), .B(n427), .ZN(n358) );
  XNOR2_X1 U425 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U426 ( .A(n360), .B(KEYINPUT14), .Z(n363) );
  XNOR2_X1 U427 ( .A(n361), .B(KEYINPUT82), .ZN(n362) );
  XNOR2_X1 U428 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n572) );
  XOR2_X1 U430 ( .A(G197GAT), .B(KEYINPUT21), .Z(n404) );
  XOR2_X1 U431 ( .A(n368), .B(n367), .Z(n370) );
  NAND2_X1 U432 ( .A1(G226GAT), .A2(G233GAT), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n372) );
  XNOR2_X1 U434 ( .A(G176GAT), .B(KEYINPUT18), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n373), .B(KEYINPUT17), .ZN(n374) );
  XOR2_X1 U436 ( .A(n374), .B(KEYINPUT19), .Z(n376) );
  XNOR2_X1 U437 ( .A(G169GAT), .B(G190GAT), .ZN(n375) );
  XOR2_X1 U438 ( .A(n376), .B(n375), .Z(n391) );
  XOR2_X1 U439 ( .A(n391), .B(n377), .Z(n378) );
  XOR2_X1 U440 ( .A(n289), .B(n378), .Z(n520) );
  XOR2_X1 U441 ( .A(G71GAT), .B(KEYINPUT20), .Z(n381) );
  XNOR2_X1 U442 ( .A(G127GAT), .B(KEYINPUT84), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n390) );
  XNOR2_X1 U444 ( .A(G113GAT), .B(KEYINPUT83), .ZN(n382) );
  XNOR2_X1 U445 ( .A(n292), .B(n382), .ZN(n428) );
  NAND2_X1 U446 ( .A1(G227GAT), .A2(G233GAT), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n293), .B(n383), .ZN(n388) );
  XNOR2_X1 U448 ( .A(G99GAT), .B(n384), .ZN(n386) );
  XNOR2_X1 U449 ( .A(n390), .B(n389), .ZN(n392) );
  XOR2_X1 U450 ( .A(G155GAT), .B(G204GAT), .Z(n394) );
  XNOR2_X1 U451 ( .A(G218GAT), .B(G211GAT), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n398) );
  XOR2_X1 U453 ( .A(KEYINPUT88), .B(KEYINPUT86), .Z(n396) );
  XNOR2_X1 U454 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n395) );
  XNOR2_X1 U455 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U456 ( .A(n398), .B(n397), .Z(n403) );
  XOR2_X1 U457 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n400) );
  NAND2_X1 U458 ( .A1(G228GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n401) );
  XNOR2_X1 U460 ( .A(G22GAT), .B(n401), .ZN(n402) );
  XNOR2_X1 U461 ( .A(n403), .B(n402), .ZN(n405) );
  XOR2_X1 U462 ( .A(n405), .B(n404), .Z(n409) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U464 ( .A(n409), .B(n408), .ZN(n413) );
  XOR2_X1 U465 ( .A(KEYINPUT2), .B(G162GAT), .Z(n411) );
  XNOR2_X1 U466 ( .A(KEYINPUT87), .B(KEYINPUT3), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U468 ( .A(G141GAT), .B(n412), .ZN(n431) );
  XNOR2_X1 U469 ( .A(n413), .B(n431), .ZN(n474) );
  NOR2_X1 U470 ( .A1(n532), .A2(n474), .ZN(n415) );
  XNOR2_X1 U471 ( .A(KEYINPUT100), .B(KEYINPUT26), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n565) );
  NAND2_X1 U473 ( .A1(n443), .A2(n565), .ZN(n420) );
  INV_X1 U474 ( .A(n520), .ZN(n470) );
  NOR2_X1 U475 ( .A1(n470), .A2(n477), .ZN(n416) );
  XNOR2_X1 U476 ( .A(KEYINPUT101), .B(n416), .ZN(n417) );
  NAND2_X1 U477 ( .A1(n417), .A2(n474), .ZN(n418) );
  XOR2_X1 U478 ( .A(KEYINPUT25), .B(n418), .Z(n419) );
  NAND2_X1 U479 ( .A1(n420), .A2(n419), .ZN(n441) );
  XOR2_X1 U480 ( .A(KEYINPUT93), .B(KEYINPUT1), .Z(n422) );
  XNOR2_X1 U481 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U483 ( .A(KEYINPUT5), .B(KEYINPUT4), .Z(n424) );
  XNOR2_X1 U484 ( .A(KEYINPUT6), .B(KEYINPUT94), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U486 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U487 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n432), .B(n431), .ZN(n440) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n438) );
  XOR2_X1 U491 ( .A(KEYINPUT92), .B(G57GAT), .Z(n434) );
  XNOR2_X1 U492 ( .A(G134GAT), .B(G148GAT), .ZN(n433) );
  XNOR2_X1 U493 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U494 ( .A(G29GAT), .B(G85GAT), .Z(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U497 ( .A(n440), .B(n439), .ZN(n442) );
  NAND2_X1 U498 ( .A1(n441), .A2(n442), .ZN(n448) );
  XNOR2_X1 U499 ( .A(KEYINPUT85), .B(n532), .ZN(n446) );
  XNOR2_X1 U500 ( .A(KEYINPUT95), .B(n442), .ZN(n517) );
  NAND2_X1 U501 ( .A1(n443), .A2(n517), .ZN(n444) );
  XOR2_X1 U502 ( .A(KEYINPUT99), .B(n444), .Z(n529) );
  NOR2_X1 U503 ( .A1(n534), .A2(n529), .ZN(n445) );
  NAND2_X1 U504 ( .A1(n446), .A2(n445), .ZN(n447) );
  NAND2_X1 U505 ( .A1(n448), .A2(n447), .ZN(n488) );
  NAND2_X1 U506 ( .A1(n572), .A2(n488), .ZN(n449) );
  XNOR2_X1 U507 ( .A(KEYINPUT106), .B(n449), .ZN(n450) );
  NOR2_X1 U508 ( .A1(n578), .A2(n450), .ZN(n452) );
  XNOR2_X1 U509 ( .A(KEYINPUT107), .B(KEYINPUT37), .ZN(n451) );
  XOR2_X1 U510 ( .A(n452), .B(n451), .Z(n515) );
  NAND2_X1 U511 ( .A1(n503), .A2(n532), .ZN(n455) );
  INV_X1 U512 ( .A(KEYINPUT123), .ZN(n480) );
  XNOR2_X1 U513 ( .A(n572), .B(KEYINPUT115), .ZN(n557) );
  XOR2_X1 U514 ( .A(n569), .B(KEYINPUT64), .Z(n456) );
  INV_X1 U515 ( .A(n546), .ZN(n457) );
  NOR2_X1 U516 ( .A1(n457), .A2(n566), .ZN(n458) );
  XNOR2_X1 U517 ( .A(n458), .B(KEYINPUT46), .ZN(n459) );
  NOR2_X1 U518 ( .A1(n557), .A2(n459), .ZN(n460) );
  INV_X1 U519 ( .A(n559), .ZN(n552) );
  AND2_X1 U520 ( .A1(n460), .A2(n552), .ZN(n462) );
  XOR2_X1 U521 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n461) );
  XNOR2_X1 U522 ( .A(n462), .B(n290), .ZN(n467) );
  NOR2_X1 U523 ( .A1(n572), .A2(n578), .ZN(n463) );
  XNOR2_X1 U524 ( .A(n463), .B(KEYINPUT45), .ZN(n464) );
  NAND2_X1 U525 ( .A1(n464), .A2(n569), .ZN(n465) );
  NOR2_X1 U526 ( .A1(n555), .A2(n465), .ZN(n466) );
  NOR2_X1 U527 ( .A1(n467), .A2(n466), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n469), .B(n468), .ZN(n530) );
  NOR2_X1 U529 ( .A1(n530), .A2(n470), .ZN(n471) );
  XNOR2_X1 U530 ( .A(n471), .B(KEYINPUT54), .ZN(n473) );
  NAND2_X1 U531 ( .A1(n294), .A2(n474), .ZN(n476) );
  XOR2_X1 U532 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n475) );
  XNOR2_X1 U533 ( .A(n476), .B(n475), .ZN(n478) );
  NOR2_X1 U534 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U535 ( .A(n480), .B(n479), .ZN(n560) );
  NAND2_X1 U536 ( .A1(n560), .A2(n546), .ZN(n483) );
  XOR2_X1 U537 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n481) );
  XNOR2_X1 U538 ( .A(n483), .B(n482), .ZN(G1349GAT) );
  NAND2_X1 U539 ( .A1(n503), .A2(n517), .ZN(n486) );
  XOR2_X1 U540 ( .A(KEYINPUT108), .B(KEYINPUT39), .Z(n484) );
  XNOR2_X1 U541 ( .A(n484), .B(G29GAT), .ZN(n485) );
  XNOR2_X1 U542 ( .A(n486), .B(n485), .ZN(G1328GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT34), .B(KEYINPUT102), .Z(n492) );
  NOR2_X1 U544 ( .A1(n572), .A2(n559), .ZN(n487) );
  XNOR2_X1 U545 ( .A(n487), .B(KEYINPUT16), .ZN(n489) );
  NAND2_X1 U546 ( .A1(n489), .A2(n488), .ZN(n507) );
  NOR2_X1 U547 ( .A1(n490), .A2(n507), .ZN(n499) );
  NAND2_X1 U548 ( .A1(n499), .A2(n517), .ZN(n491) );
  XNOR2_X1 U549 ( .A(n492), .B(n491), .ZN(n493) );
  XOR2_X1 U550 ( .A(G1GAT), .B(n493), .Z(G1324GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n495) );
  NAND2_X1 U552 ( .A1(n499), .A2(n520), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U554 ( .A(G8GAT), .B(n496), .ZN(G1325GAT) );
  XOR2_X1 U555 ( .A(G15GAT), .B(KEYINPUT35), .Z(n498) );
  NAND2_X1 U556 ( .A1(n499), .A2(n532), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(G1326GAT) );
  XOR2_X1 U558 ( .A(G22GAT), .B(KEYINPUT105), .Z(n501) );
  NAND2_X1 U559 ( .A1(n499), .A2(n534), .ZN(n500) );
  XNOR2_X1 U560 ( .A(n501), .B(n500), .ZN(G1327GAT) );
  NAND2_X1 U561 ( .A1(n520), .A2(n503), .ZN(n502) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n502), .ZN(G1329GAT) );
  XOR2_X1 U563 ( .A(G50GAT), .B(KEYINPUT109), .Z(n505) );
  NAND2_X1 U564 ( .A1(n534), .A2(n503), .ZN(n504) );
  XNOR2_X1 U565 ( .A(n505), .B(n504), .ZN(G1331GAT) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n509) );
  NAND2_X1 U567 ( .A1(n546), .A2(n566), .ZN(n506) );
  XNOR2_X1 U568 ( .A(n506), .B(KEYINPUT110), .ZN(n516) );
  NOR2_X1 U569 ( .A1(n516), .A2(n507), .ZN(n512) );
  NAND2_X1 U570 ( .A1(n512), .A2(n517), .ZN(n508) );
  XNOR2_X1 U571 ( .A(n509), .B(n508), .ZN(G1332GAT) );
  NAND2_X1 U572 ( .A1(n520), .A2(n512), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n510), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U574 ( .A1(n512), .A2(n532), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U576 ( .A(G78GAT), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U577 ( .A1(n512), .A2(n534), .ZN(n513) );
  XNOR2_X1 U578 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  XOR2_X1 U579 ( .A(G85GAT), .B(KEYINPUT111), .Z(n519) );
  NOR2_X1 U580 ( .A1(n516), .A2(n515), .ZN(n524) );
  NAND2_X1 U581 ( .A1(n524), .A2(n517), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n519), .B(n518), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n520), .A2(n524), .ZN(n521) );
  XNOR2_X1 U584 ( .A(n521), .B(KEYINPUT112), .ZN(n522) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n522), .ZN(G1337GAT) );
  NAND2_X1 U586 ( .A1(n524), .A2(n532), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n528) );
  XOR2_X1 U589 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n526) );
  NAND2_X1 U590 ( .A1(n524), .A2(n534), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n528), .B(n527), .ZN(G1339GAT) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(KEYINPUT120), .ZN(n536) );
  NOR2_X1 U594 ( .A1(n530), .A2(n529), .ZN(n531) );
  XOR2_X1 U595 ( .A(KEYINPUT119), .B(n531), .Z(n544) );
  NAND2_X1 U596 ( .A1(n532), .A2(n544), .ZN(n533) );
  NOR2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n541), .A2(n555), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n536), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U601 ( .A1(n541), .A2(n546), .ZN(n537) );
  XNOR2_X1 U602 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  NAND2_X1 U603 ( .A1(n557), .A2(n541), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n539), .B(KEYINPUT50), .ZN(n540) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U607 ( .A1(n541), .A2(n559), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(G1343GAT) );
  NAND2_X1 U609 ( .A1(n565), .A2(n544), .ZN(n551) );
  NOR2_X1 U610 ( .A1(n566), .A2(n551), .ZN(n545) );
  XOR2_X1 U611 ( .A(G141GAT), .B(n545), .Z(G1344GAT) );
  NOR2_X1 U612 ( .A1(n457), .A2(n551), .ZN(n548) );
  XNOR2_X1 U613 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G148GAT), .B(n549), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n572), .A2(n551), .ZN(n550) );
  XOR2_X1 U617 ( .A(G155GAT), .B(n550), .Z(G1346GAT) );
  NOR2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(KEYINPUT121), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n560), .A2(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n557), .A2(n560), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U625 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n562) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1351GAT) );
  XOR2_X1 U628 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n564) );
  XNOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n568) );
  NAND2_X1 U631 ( .A1(n294), .A2(n565), .ZN(n577) );
  NOR2_X1 U632 ( .A1(n566), .A2(n577), .ZN(n567) );
  XOR2_X1 U633 ( .A(n568), .B(n567), .Z(G1352GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n577), .ZN(n571) );
  XNOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n577), .ZN(n574) );
  XNOR2_X1 U638 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(G1354GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n576) );
  XNOR2_X1 U641 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(n580) );
  NOR2_X1 U643 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U644 ( .A(n580), .B(n579), .Z(G1355GAT) );
endmodule

