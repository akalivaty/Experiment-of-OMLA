//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 0 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n613, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  INV_X1    g022(.A(G567), .ZN(new_n448));
  NOR2_X1   g023(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT64), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  OAI21_X1  g033(.A(new_n458), .B1(new_n448), .B2(new_n454), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT65), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  OR2_X1    g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n471), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n468), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  NOR2_X1   g051(.A1(new_n465), .A2(new_n472), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n477), .A2(G124), .B1(G136), .B2(new_n471), .ZN(new_n478));
  INV_X1    g053(.A(G100), .ZN(new_n479));
  AND3_X1   g054(.A1(new_n479), .A2(new_n472), .A3(KEYINPUT66), .ZN(new_n480));
  AOI21_X1  g055(.A(KEYINPUT66), .B1(new_n479), .B2(new_n472), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G112), .B2(new_n472), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n478), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g058(.A(new_n483), .B(KEYINPUT67), .Z(G162));
  OAI21_X1  g059(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n485), .B1(new_n486), .B2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n469), .A2(new_n470), .ZN(new_n489));
  AND2_X1   g064(.A1(G126), .A2(G2105), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT68), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(KEYINPUT68), .B(new_n490), .C1(new_n463), .C2(new_n464), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n488), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n490), .B1(new_n463), .B2(new_n464), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n487), .B1(new_n499), .B2(new_n492), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT69), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n472), .C1(new_n463), .C2(new_n464), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT4), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n489), .A2(new_n504), .A3(G138), .A4(new_n472), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n496), .A2(new_n501), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n509), .A2(G62), .ZN(new_n510));
  NAND2_X1  g085(.A1(G75), .A2(G543), .ZN(new_n511));
  XOR2_X1   g086(.A(new_n511), .B(KEYINPUT71), .Z(new_n512));
  OAI21_X1  g087(.A(G651), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT72), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT70), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(G651), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  OAI21_X1  g097(.A(new_n515), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G543), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n524), .B1(new_n518), .B2(new_n519), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n525), .A2(KEYINPUT70), .A3(G50), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n520), .A2(new_n509), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n523), .A2(new_n526), .B1(G88), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT72), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n529), .B(G651), .C1(new_n510), .C2(new_n512), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n514), .A2(new_n528), .A3(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  NAND2_X1  g107(.A1(new_n525), .A2(G51), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n520), .A2(new_n509), .ZN(new_n534));
  XOR2_X1   g109(.A(KEYINPUT73), .B(G89), .Z(new_n535));
  OAI21_X1  g110(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n536), .A2(new_n540), .ZN(G168));
  NAND2_X1  g116(.A1(new_n525), .A2(G52), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n534), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n517), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n544), .A2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n525), .A2(G43), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n549), .B2(new_n534), .ZN(new_n550));
  AOI22_X1  g125(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n517), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  NAND4_X1  g129(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND4_X1  g132(.A1(G319), .A2(G483), .A3(G661), .A4(new_n557), .ZN(G188));
  AOI22_X1  g133(.A1(new_n509), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n559));
  OR2_X1    g134(.A1(new_n559), .A2(new_n517), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n527), .A2(G91), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OAI211_X1 g138(.A(KEYINPUT74), .B(new_n562), .C1(new_n521), .C2(new_n563), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT74), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n563), .B1(new_n565), .B2(KEYINPUT9), .ZN(new_n566));
  OAI211_X1 g141(.A(new_n525), .B(new_n566), .C1(new_n565), .C2(KEYINPUT9), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n560), .A2(new_n561), .A3(new_n564), .A4(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  NAND2_X1  g145(.A1(new_n527), .A2(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n525), .A2(G49), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(G73), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(new_n509), .ZN(new_n576));
  INV_X1    g151(.A(G61), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n578), .A2(G651), .B1(G48), .B2(new_n525), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n520), .A2(new_n509), .A3(G86), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT75), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n520), .A2(new_n509), .A3(KEYINPUT75), .A4(G86), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n579), .A2(new_n584), .ZN(G305));
  NAND2_X1  g160(.A1(new_n525), .A2(G47), .ZN(new_n586));
  XNOR2_X1  g161(.A(KEYINPUT76), .B(G85), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n534), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(KEYINPUT77), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n586), .B(new_n590), .C1(new_n534), .C2(new_n587), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n509), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n517), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n592), .A2(new_n594), .ZN(G290));
  NAND3_X1  g170(.A1(new_n527), .A2(KEYINPUT10), .A3(G92), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT10), .ZN(new_n597));
  INV_X1    g172(.A(G92), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n534), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n576), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n603), .A2(G651), .B1(G54), .B2(new_n525), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n607), .B1(new_n606), .B2(G171), .ZN(G284));
  OAI21_X1  g183(.A(new_n607), .B1(new_n606), .B2(G171), .ZN(G321));
  NAND2_X1  g184(.A1(G299), .A2(new_n606), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(new_n606), .B2(G168), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(new_n606), .B2(G168), .ZN(G280));
  AND2_X1   g187(.A1(new_n600), .A2(new_n604), .ZN(new_n613));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n613), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n489), .A2(new_n473), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT12), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT12), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n489), .A2(new_n622), .A3(new_n473), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  INV_X1    g200(.A(G2100), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n477), .A2(G123), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n471), .A2(G135), .ZN(new_n630));
  NOR2_X1   g205(.A1(new_n472), .A2(G111), .ZN(new_n631));
  OAI21_X1  g206(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n629), .B(new_n630), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(G2096), .Z(new_n634));
  NAND3_X1  g209(.A1(new_n627), .A2(new_n628), .A3(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(G1341), .B(G1348), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2427), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2430), .ZN(new_n638));
  XNOR2_X1  g213(.A(KEYINPUT15), .B(G2435), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2451), .B(G2454), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT16), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2443), .B(G2446), .ZN(new_n646));
  INV_X1    g221(.A(new_n644), .ZN(new_n647));
  NAND4_X1  g222(.A1(new_n640), .A2(KEYINPUT14), .A3(new_n647), .A4(new_n641), .ZN(new_n648));
  AND3_X1   g223(.A1(new_n645), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n646), .B1(new_n645), .B2(new_n648), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n636), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT78), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n649), .A2(new_n650), .A3(new_n636), .ZN(new_n654));
  INV_X1    g229(.A(G14), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n653), .A2(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2084), .B(G2090), .Z(new_n658));
  XNOR2_X1  g233(.A(G2067), .B(G2678), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G2072), .B(G2078), .Z(new_n661));
  NOR2_X1   g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n661), .B(KEYINPUT17), .ZN(new_n664));
  INV_X1    g239(.A(new_n658), .ZN(new_n665));
  INV_X1    g240(.A(new_n659), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n665), .A2(new_n661), .A3(new_n666), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(new_n660), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n663), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2096), .B(G2100), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT79), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n670), .B(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1991), .B(G1996), .Z(new_n674));
  XOR2_X1   g249(.A(KEYINPUT80), .B(KEYINPUT19), .Z(new_n675));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n678), .A2(KEYINPUT81), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(KEYINPUT81), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  OR3_X1    g258(.A1(new_n677), .A2(new_n683), .A3(KEYINPUT20), .ZN(new_n684));
  OAI21_X1  g259(.A(KEYINPUT20), .B1(new_n677), .B2(new_n683), .ZN(new_n685));
  AND2_X1   g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(KEYINPUT82), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n678), .B(KEYINPUT81), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n688), .A2(new_n681), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n689), .A2(new_n677), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n689), .A2(new_n683), .A3(new_n677), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n686), .A2(new_n687), .A3(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n690), .A2(new_n691), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n684), .A2(new_n685), .ZN(new_n695));
  AOI21_X1  g270(.A(KEYINPUT82), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g273(.A1(new_n693), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n687), .B1(new_n686), .B2(new_n692), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n694), .A2(new_n695), .A3(KEYINPUT82), .ZN(new_n701));
  AOI21_X1  g276(.A(new_n697), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n674), .B1(new_n699), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1981), .B(G1986), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n698), .B1(new_n693), .B2(new_n696), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n700), .A2(new_n701), .A3(new_n697), .ZN(new_n706));
  INV_X1    g281(.A(new_n674), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n705), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n703), .A2(new_n704), .A3(new_n708), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n704), .B1(new_n703), .B2(new_n708), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(G229));
  NAND2_X1  g286(.A1(new_n477), .A2(G119), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n471), .A2(G131), .ZN(new_n713));
  OR2_X1    g288(.A1(G95), .A2(G2105), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n714), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  MUX2_X1   g291(.A(G25), .B(new_n716), .S(G29), .Z(new_n717));
  XOR2_X1   g292(.A(KEYINPUT35), .B(G1991), .Z(new_n718));
  INV_X1    g293(.A(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n717), .B(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G24), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT83), .ZN(new_n723));
  INV_X1    g298(.A(G290), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n721), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(G1986), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n721), .A2(G6), .ZN(new_n727));
  INV_X1    g302(.A(G305), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n727), .B1(new_n728), .B2(new_n721), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT84), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT32), .B(G1981), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n721), .A2(G23), .ZN(new_n733));
  INV_X1    g308(.A(G288), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(new_n721), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT85), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT33), .B(G1976), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n736), .B(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(G16), .A2(G22), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G166), .B2(G16), .ZN(new_n740));
  INV_X1    g315(.A(G1971), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n732), .A2(new_n738), .A3(new_n742), .ZN(new_n743));
  AOI211_X1 g318(.A(new_n720), .B(new_n726), .C1(new_n743), .C2(KEYINPUT34), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(KEYINPUT34), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT36), .ZN(new_n747));
  INV_X1    g322(.A(G29), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n748), .A2(G35), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G162), .B2(new_n748), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT29), .Z(new_n751));
  INV_X1    g326(.A(G2090), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT93), .B(KEYINPUT24), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G34), .ZN(new_n755));
  MUX2_X1   g330(.A(new_n755), .B(new_n475), .S(G29), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n756), .A2(G2084), .ZN(new_n757));
  NOR2_X1   g332(.A1(G171), .A2(new_n721), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G5), .B2(new_n721), .ZN(new_n759));
  INV_X1    g334(.A(G1961), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G168), .A2(new_n721), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n721), .B2(G21), .ZN(new_n763));
  INV_X1    g338(.A(G1966), .ZN(new_n764));
  OAI22_X1  g339(.A1(new_n763), .A2(new_n764), .B1(new_n756), .B2(G2084), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT30), .B(G28), .ZN(new_n767));
  OR2_X1    g342(.A1(KEYINPUT31), .A2(G11), .ZN(new_n768));
  NAND2_X1  g343(.A1(KEYINPUT31), .A2(G11), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n767), .A2(new_n748), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n633), .B2(new_n748), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n763), .B2(new_n764), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n748), .A2(G32), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n477), .A2(G129), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n471), .A2(G141), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n473), .A2(G105), .ZN(new_n776));
  AND3_X1   g351(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT94), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT26), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n773), .B1(new_n782), .B2(new_n748), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT27), .B(G1996), .Z(new_n784));
  OAI211_X1 g359(.A(new_n766), .B(new_n772), .C1(new_n783), .C2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(G4), .A2(G16), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n613), .B2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT86), .B(G1348), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(G115), .A2(G2104), .ZN(new_n790));
  INV_X1    g365(.A(G127), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n465), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n792), .A2(G2105), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT25), .ZN(new_n794));
  NAND2_X1  g369(.A1(G103), .A2(G2104), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(G2105), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n472), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n471), .A2(G139), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(new_n748), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n748), .B2(G33), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT92), .B(G2072), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n759), .A2(new_n760), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n802), .A2(new_n803), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n789), .A2(new_n804), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NOR3_X1   g382(.A1(new_n753), .A2(new_n785), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(new_n751), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n808), .B1(G2090), .B2(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(G104), .A2(G2105), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n811), .B(G2104), .C1(G116), .C2(new_n472), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT88), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n477), .A2(G128), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n471), .A2(G140), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(KEYINPUT89), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(KEYINPUT88), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n812), .B(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(KEYINPUT89), .ZN(new_n820));
  NAND4_X1  g395(.A1(new_n819), .A2(new_n820), .A3(new_n815), .A4(new_n814), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(G29), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(KEYINPUT90), .ZN(new_n824));
  XOR2_X1   g399(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n825));
  NAND2_X1  g400(.A1(new_n748), .A2(G26), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G2067), .ZN(new_n829));
  NOR2_X1   g404(.A1(G164), .A2(new_n748), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(G27), .B2(new_n748), .ZN(new_n831));
  INV_X1    g406(.A(G2078), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g408(.A(G19), .ZN(new_n834));
  OR3_X1    g409(.A1(new_n834), .A2(KEYINPUT87), .A3(G16), .ZN(new_n835));
  OAI21_X1  g410(.A(KEYINPUT87), .B1(new_n834), .B2(G16), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n835), .B(new_n836), .C1(new_n553), .C2(new_n721), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G1341), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n721), .A2(G20), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT95), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT23), .ZN(new_n841));
  INV_X1    g416(.A(G299), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n841), .B1(new_n842), .B2(new_n721), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT96), .B(G1956), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n838), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n831), .A2(new_n832), .ZN(new_n847));
  INV_X1    g422(.A(new_n843), .ZN(new_n848));
  AOI22_X1  g423(.A1(new_n848), .A2(new_n844), .B1(new_n783), .B2(new_n784), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  NOR4_X1   g425(.A1(new_n810), .A2(new_n829), .A3(new_n833), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n747), .A2(new_n851), .ZN(G150));
  INV_X1    g427(.A(G150), .ZN(G311));
  INV_X1    g428(.A(G93), .ZN(new_n854));
  XOR2_X1   g429(.A(KEYINPUT97), .B(G55), .Z(new_n855));
  OAI22_X1  g430(.A1(new_n854), .A2(new_n534), .B1(new_n521), .B2(new_n855), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n509), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(new_n517), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT99), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  OAI21_X1  g436(.A(KEYINPUT99), .B1(new_n856), .B2(new_n858), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(G860), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(KEYINPUT37), .Z(new_n865));
  NAND2_X1  g440(.A1(new_n613), .A2(G559), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT38), .ZN(new_n867));
  OR2_X1    g442(.A1(new_n550), .A2(new_n552), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n861), .A2(new_n868), .A3(new_n862), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n553), .B(KEYINPUT98), .C1(new_n858), .C2(new_n856), .ZN(new_n870));
  INV_X1    g445(.A(KEYINPUT98), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n868), .B2(new_n859), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n869), .A2(new_n870), .A3(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n867), .B(new_n873), .Z(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n875), .A2(KEYINPUT39), .ZN(new_n876));
  INV_X1    g451(.A(G860), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(new_n875), .B2(KEYINPUT39), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n865), .B1(new_n876), .B2(new_n878), .ZN(G145));
  AOI21_X1  g454(.A(new_n504), .B1(new_n471), .B2(G138), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n881));
  OAI21_X1  g456(.A(KEYINPUT100), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n503), .A2(new_n505), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n500), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n822), .A2(new_n885), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n882), .A2(new_n500), .A3(new_n884), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(new_n817), .A3(new_n821), .ZN(new_n888));
  OAI21_X1  g463(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n889));
  INV_X1    g464(.A(G118), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n889), .B1(new_n890), .B2(G2105), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n891), .B1(new_n477), .B2(G130), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n471), .A2(KEYINPUT101), .A3(G142), .ZN(new_n893));
  AOI21_X1  g468(.A(KEYINPUT101), .B1(new_n471), .B2(G142), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n886), .A2(new_n888), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n895), .B1(new_n886), .B2(new_n888), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n781), .A2(new_n799), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n800), .A2(new_n777), .A3(new_n780), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n716), .A2(new_n621), .A3(new_n623), .ZN(new_n901));
  NAND4_X1  g476(.A1(new_n624), .A2(new_n713), .A3(new_n712), .A4(new_n715), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AND3_X1   g478(.A1(new_n899), .A2(new_n900), .A3(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n903), .B1(new_n899), .B2(new_n900), .ZN(new_n905));
  OAI22_X1  g480(.A1(new_n897), .A2(new_n898), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n904), .A2(new_n905), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n886), .A2(new_n888), .ZN(new_n908));
  INV_X1    g483(.A(new_n895), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n907), .A2(new_n910), .A3(new_n896), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n906), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(G160), .A2(new_n633), .ZN(new_n913));
  OR2_X1    g488(.A1(G160), .A2(new_n633), .ZN(new_n914));
  NAND3_X1  g489(.A1(G162), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT103), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n913), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n483), .B(KEYINPUT67), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n915), .A2(new_n916), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n916), .B1(new_n915), .B2(new_n919), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n912), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(G37), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n906), .A2(new_n911), .A3(new_n915), .A4(new_n919), .ZN(new_n926));
  OR2_X1    g501(.A1(new_n926), .A2(KEYINPUT102), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(KEYINPUT102), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g504(.A(KEYINPUT104), .B(KEYINPUT40), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n929), .B(new_n930), .ZN(G395));
  XOR2_X1   g506(.A(new_n873), .B(new_n616), .Z(new_n932));
  NAND2_X1  g507(.A1(new_n842), .A2(new_n605), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT105), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n613), .A2(G299), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n842), .A2(new_n936), .A3(new_n605), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n934), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n939), .B1(new_n613), .B2(G299), .ZN(new_n940));
  AOI22_X1  g515(.A1(new_n938), .A2(new_n939), .B1(new_n933), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n942));
  OR3_X1    g517(.A1(new_n932), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n933), .A2(new_n935), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n932), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n942), .B1(new_n932), .B2(new_n941), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n947), .B(KEYINPUT42), .Z(new_n948));
  XNOR2_X1  g523(.A(G305), .B(KEYINPUT108), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(G303), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n728), .A2(KEYINPUT108), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n579), .A2(KEYINPUT108), .A3(new_n584), .ZN(new_n952));
  OAI21_X1  g527(.A(G166), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(G290), .A2(KEYINPUT107), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT107), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n592), .A2(new_n956), .A3(new_n594), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n957), .A3(new_n734), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n955), .A2(new_n957), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(G288), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n954), .A2(KEYINPUT109), .A3(new_n958), .A4(new_n960), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(KEYINPUT109), .A3(new_n958), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n950), .A2(new_n953), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT109), .B1(new_n960), .B2(new_n958), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n948), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n948), .A2(new_n967), .ZN(new_n969));
  OAI21_X1  g544(.A(G868), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n863), .A2(new_n606), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(G295));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n971), .ZN(G331));
  XNOR2_X1  g548(.A(G171), .B(G168), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n974), .A2(new_n869), .A3(new_n870), .A4(new_n872), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n975), .A2(new_n944), .ZN(new_n976));
  INV_X1    g551(.A(new_n974), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n873), .A2(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT110), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n873), .A2(new_n977), .A3(KEYINPUT110), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n976), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n978), .A2(new_n975), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n982), .B1(new_n941), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n924), .B1(new_n966), .B2(new_n984), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n941), .A2(new_n983), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n960), .A2(new_n958), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT109), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(new_n962), .A3(new_n963), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n986), .A2(new_n982), .B1(new_n990), .B2(new_n961), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT43), .B1(new_n985), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n976), .A2(new_n978), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n980), .A2(new_n975), .A3(new_n981), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n934), .A2(new_n937), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n995), .A2(new_n940), .B1(new_n939), .B2(new_n944), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n993), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(new_n966), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n986), .A2(new_n990), .A3(new_n961), .A4(new_n982), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n998), .A2(new_n999), .A3(new_n1000), .A4(new_n924), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n992), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1002), .A2(KEYINPUT44), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n985), .B1(new_n966), .B2(new_n997), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT111), .ZN(new_n1005));
  OR3_X1    g580(.A1(new_n1004), .A2(new_n1005), .A3(new_n1000), .ZN(new_n1006));
  OR3_X1    g581(.A1(new_n985), .A2(new_n991), .A3(KEYINPUT43), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n1005), .B1(new_n1004), .B2(new_n1000), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1003), .B1(new_n1009), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n885), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AND3_X1   g589(.A1(new_n468), .A2(G40), .A3(new_n474), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G2067), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n822), .B(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1018), .B1(new_n1020), .B2(new_n782), .ZN(new_n1021));
  INV_X1    g596(.A(G1996), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1017), .A2(KEYINPUT46), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT46), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1024));
  NOR3_X1   g599(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  XOR2_X1   g600(.A(new_n1025), .B(KEYINPUT47), .Z(new_n1026));
  XNOR2_X1  g601(.A(new_n781), .B(new_n1022), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1020), .A2(new_n1027), .ZN(new_n1028));
  OR2_X1    g603(.A1(new_n716), .A2(new_n719), .ZN(new_n1029));
  OAI22_X1  g604(.A1(new_n1028), .A2(new_n1029), .B1(G2067), .B2(new_n822), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1030), .A2(new_n1017), .ZN(new_n1031));
  XOR2_X1   g606(.A(new_n1031), .B(KEYINPUT125), .Z(new_n1032));
  NAND2_X1  g607(.A1(new_n716), .A2(new_n719), .ZN(new_n1033));
  AND4_X1   g608(.A1(new_n1020), .A2(new_n1027), .A3(new_n1029), .A4(new_n1033), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(new_n1018), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT48), .ZN(new_n1036));
  OR3_X1    g611(.A1(new_n1018), .A2(G1986), .A3(G290), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1038), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1039));
  AND3_X1   g614(.A1(new_n1026), .A2(new_n1032), .A3(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n885), .A2(new_n1011), .A3(new_n1015), .ZN(new_n1041));
  INV_X1    g616(.A(G1981), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n579), .A2(new_n1042), .A3(new_n584), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n525), .A2(G48), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n509), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n1045));
  OAI211_X1 g620(.A(new_n1044), .B(new_n580), .C1(new_n1045), .C2(new_n517), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G1981), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT49), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1043), .A2(KEYINPUT49), .A3(new_n1047), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1050), .A2(G8), .A3(new_n1041), .A4(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1052), .A2(new_n1053), .A3(new_n734), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1043), .ZN(new_n1055));
  OAI211_X1 g630(.A(G8), .B(new_n1041), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n885), .A2(KEYINPUT45), .A3(new_n1011), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n1015), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT45), .B1(new_n507), .B2(new_n1011), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n741), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n506), .B1(new_n500), .B2(KEYINPUT69), .ZN(new_n1061));
  AOI211_X1 g636(.A(new_n495), .B(new_n487), .C1(new_n499), .C2(new_n492), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1011), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT50), .ZN(new_n1064));
  XNOR2_X1  g639(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n885), .A2(new_n1011), .A3(new_n1065), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1064), .A2(new_n752), .A3(new_n1015), .A4(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1060), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(G303), .A2(G8), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT55), .ZN(new_n1070));
  XNOR2_X1  g645(.A(new_n1069), .B(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1068), .A2(G8), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n734), .A2(G1976), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1041), .A2(new_n1073), .A3(G8), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(KEYINPUT52), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1041), .A2(new_n1073), .A3(G8), .A4(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1052), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1056), .B1(new_n1072), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1078), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1072), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT63), .ZN(new_n1082));
  INV_X1    g657(.A(G8), .ZN(new_n1083));
  OAI211_X1 g658(.A(KEYINPUT45), .B(new_n1011), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n883), .B1(new_n503), .B2(new_n505), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1085), .A2(new_n494), .ZN(new_n1086));
  AOI21_X1  g661(.A(G1384), .B1(new_n1086), .B2(new_n884), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1084), .B(new_n1015), .C1(new_n1087), .C2(KEYINPUT45), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n764), .ZN(new_n1089));
  INV_X1    g664(.A(G2084), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1064), .A2(new_n1090), .A3(new_n1015), .A4(new_n1066), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1083), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(G168), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1081), .A2(new_n1082), .A3(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1083), .B1(new_n1060), .B2(new_n1067), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1095), .A2(KEYINPUT113), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1071), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1095), .B2(KEYINPUT113), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1094), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1065), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1012), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT50), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n507), .A2(new_n1102), .A3(new_n1011), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(new_n1103), .A3(new_n1015), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1060), .B1(G2090), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(G8), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n1097), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1078), .B1(new_n1095), .B2(new_n1071), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1082), .B1(new_n1109), .B2(new_n1093), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1079), .B1(new_n1099), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1089), .A2(G168), .A3(new_n1091), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(G8), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT51), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(KEYINPUT51), .A3(G8), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(KEYINPUT120), .A3(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT51), .B1(new_n1112), .B2(G8), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  AOI22_X1  g694(.A1(new_n1118), .A2(new_n1119), .B1(G286), .B2(new_n1092), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT62), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1117), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1063), .A2(new_n1013), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1125), .A2(new_n832), .A3(new_n1015), .A4(new_n1057), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT53), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1066), .A2(new_n1015), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1102), .B1(new_n507), .B2(new_n1011), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n760), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1127), .A2(G2078), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1014), .A2(new_n1015), .A3(new_n1084), .A4(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1128), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(G171), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT121), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1134), .A2(new_n1137), .A3(G171), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT123), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1071), .B1(new_n1105), .B2(G8), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n1081), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1107), .A2(new_n1108), .A3(KEYINPUT123), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1124), .A2(new_n1139), .A3(new_n1142), .A4(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1111), .B1(new_n1123), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT122), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT53), .B1(new_n1146), .B2(new_n832), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1147), .B1(new_n1146), .B2(new_n832), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1014), .A2(new_n1015), .A3(new_n1057), .A4(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1128), .A2(new_n1131), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(G171), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1128), .A2(new_n1131), .A3(G301), .A4(new_n1133), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(KEYINPUT54), .A3(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1142), .A2(new_n1143), .A3(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1121), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1150), .A2(G171), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1156), .B1(new_n1139), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(KEYINPUT124), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  AND3_X1   g734(.A1(new_n1142), .A2(new_n1143), .A3(new_n1153), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1161));
  AND4_X1   g736(.A1(KEYINPUT124), .A2(new_n1160), .A3(new_n1158), .A4(new_n1161), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1159), .A2(new_n1162), .ZN(new_n1163));
  XNOR2_X1  g738(.A(KEYINPUT56), .B(G2072), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1125), .A2(new_n1015), .A3(new_n1057), .A4(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT115), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(G1956), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1104), .A2(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1016), .B1(new_n1087), .B2(KEYINPUT45), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1170), .A2(KEYINPUT115), .A3(new_n1125), .A4(new_n1164), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT114), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT57), .ZN(new_n1173));
  OAI21_X1  g748(.A(G299), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1167), .A2(new_n1169), .A3(new_n1171), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT116), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT61), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  OR2_X1    g754(.A1(new_n1179), .A2(KEYINPUT117), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1170), .A2(new_n1022), .A3(new_n1125), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1041), .ZN(new_n1182));
  XNOR2_X1  g757(.A(KEYINPUT58), .B(G1341), .ZN(new_n1183));
  OAI21_X1  g758(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(new_n553), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT59), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1177), .A2(KEYINPUT61), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1184), .A2(KEYINPUT59), .A3(new_n553), .ZN(new_n1189));
  AND3_X1   g764(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1179), .A2(KEYINPUT117), .ZN(new_n1191));
  INV_X1    g766(.A(G1348), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1192), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1193));
  NAND3_X1  g768(.A1(new_n1087), .A2(new_n1019), .A3(new_n1015), .ZN(new_n1194));
  AND2_X1   g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1195), .A2(KEYINPUT60), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1193), .A2(KEYINPUT60), .A3(new_n1194), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT118), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1197), .A2(new_n1198), .A3(new_n605), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1200), .A2(new_n613), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1202));
  OAI211_X1 g777(.A(new_n1196), .B(new_n1199), .C1(new_n1201), .C2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g778(.A1(new_n1180), .A2(new_n1190), .A3(new_n1191), .A4(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(KEYINPUT119), .ZN(new_n1205));
  AND2_X1   g780(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1176), .B1(new_n1206), .B2(new_n1171), .ZN(new_n1207));
  NOR2_X1   g782(.A1(new_n1195), .A2(new_n605), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1177), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  AND3_X1   g784(.A1(new_n1204), .A2(new_n1205), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1205), .B1(new_n1204), .B2(new_n1209), .ZN(new_n1211));
  NOR2_X1   g786(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1145), .B1(new_n1163), .B2(new_n1212), .ZN(new_n1213));
  XOR2_X1   g788(.A(G290), .B(G1986), .Z(new_n1214));
  AOI21_X1  g789(.A(new_n1018), .B1(new_n1034), .B2(new_n1214), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1040), .B1(new_n1213), .B2(new_n1215), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n1218));
  OR2_X1    g792(.A1(new_n460), .A2(G227), .ZN(new_n1219));
  AOI21_X1  g793(.A(new_n1219), .B1(new_n653), .B2(new_n656), .ZN(new_n1220));
  OAI21_X1  g794(.A(new_n1220), .B1(new_n709), .B2(new_n710), .ZN(new_n1221));
  NOR2_X1   g795(.A1(new_n929), .A2(new_n1221), .ZN(new_n1222));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n1223));
  AND3_X1   g797(.A1(new_n1002), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1224));
  AOI21_X1  g798(.A(new_n1223), .B1(new_n1002), .B2(new_n1222), .ZN(new_n1225));
  OAI21_X1  g799(.A(new_n1218), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g800(.A1(new_n1002), .A2(new_n1222), .ZN(new_n1227));
  NAND2_X1  g801(.A1(new_n1227), .A2(KEYINPUT126), .ZN(new_n1228));
  NAND3_X1  g802(.A1(new_n1002), .A2(new_n1222), .A3(new_n1223), .ZN(new_n1229));
  NAND3_X1  g803(.A1(new_n1228), .A2(KEYINPUT127), .A3(new_n1229), .ZN(new_n1230));
  AND2_X1   g804(.A1(new_n1226), .A2(new_n1230), .ZN(G308));
  NAND2_X1  g805(.A1(new_n1228), .A2(new_n1229), .ZN(G225));
endmodule


