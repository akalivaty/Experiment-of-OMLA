

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757;

  AND2_X1 U363 ( .A1(n430), .A2(n447), .ZN(n411) );
  XNOR2_X1 U364 ( .A(n743), .B(n499), .ZN(n397) );
  XOR2_X1 U365 ( .A(G902), .B(KEYINPUT15), .Z(n529) );
  INV_X1 U366 ( .A(G143), .ZN(n419) );
  AND2_X1 U367 ( .A1(n442), .A2(n412), .ZN(n341) );
  XOR2_X2 U368 ( .A(KEYINPUT45), .B(KEYINPUT85), .Z(n595) );
  NAND2_X1 U369 ( .A1(n341), .A2(n413), .ZN(n446) );
  XOR2_X1 U370 ( .A(G143), .B(G104), .Z(n545) );
  XNOR2_X2 U371 ( .A(n525), .B(G134), .ZN(n398) );
  XNOR2_X2 U372 ( .A(n580), .B(n579), .ZN(n683) );
  INV_X1 U373 ( .A(G472), .ZN(n377) );
  NOR2_X1 U374 ( .A1(n712), .A2(n381), .ZN(n713) );
  XNOR2_X1 U375 ( .A(n431), .B(n595), .ZN(n705) );
  AND2_X2 U376 ( .A1(n420), .A2(n495), .ZN(n746) );
  XNOR2_X1 U377 ( .A(n367), .B(KEYINPUT35), .ZN(n755) );
  XNOR2_X1 U378 ( .A(n625), .B(n448), .ZN(n756) );
  NOR2_X1 U379 ( .A1(n624), .A2(n635), .ZN(n625) );
  XNOR2_X1 U380 ( .A(n454), .B(KEYINPUT39), .ZN(n635) );
  AND2_X1 U381 ( .A1(n392), .A2(n390), .ZN(n454) );
  AND2_X1 U382 ( .A1(n613), .A2(n391), .ZN(n390) );
  INV_X1 U383 ( .A(n690), .ZN(n575) );
  XNOR2_X1 U384 ( .A(n383), .B(n382), .ZN(n588) );
  XNOR2_X1 U385 ( .A(n558), .B(n557), .ZN(n589) );
  OR2_X1 U386 ( .A1(n727), .A2(G902), .ZN(n439) );
  XNOR2_X1 U387 ( .A(n459), .B(n458), .ZN(n561) );
  XOR2_X1 U388 ( .A(G125), .B(G146), .Z(n523) );
  XNOR2_X2 U389 ( .A(n342), .B(n343), .ZN(n689) );
  NOR2_X1 U390 ( .A1(n573), .A2(G902), .ZN(n342) );
  XNOR2_X1 U391 ( .A(KEYINPUT100), .B(G472), .ZN(n343) );
  NOR2_X1 U392 ( .A1(n604), .A2(n542), .ZN(n423) );
  XNOR2_X1 U393 ( .A(n441), .B(n534), .ZN(n604) );
  NOR2_X1 U394 ( .A1(n474), .A2(n479), .ZN(n344) );
  INV_X1 U395 ( .A(n546), .ZN(n497) );
  XNOR2_X1 U396 ( .A(n398), .B(n497), .ZN(n385) );
  XNOR2_X1 U397 ( .A(n385), .B(n498), .ZN(n743) );
  BUF_X1 U398 ( .A(n581), .Z(n345) );
  XNOR2_X1 U399 ( .A(n423), .B(n543), .ZN(n581) );
  NAND2_X1 U400 ( .A1(n748), .A2(G224), .ZN(n417) );
  INV_X1 U401 ( .A(KEYINPUT44), .ZN(n433) );
  INV_X1 U402 ( .A(KEYINPUT8), .ZN(n458) );
  NAND2_X1 U403 ( .A1(n451), .A2(G234), .ZN(n459) );
  NAND2_X1 U404 ( .A1(n388), .A2(n461), .ZN(n387) );
  XNOR2_X1 U405 ( .A(n389), .B(n358), .ZN(n388) );
  XNOR2_X1 U406 ( .A(G113), .B(G122), .ZN(n544) );
  AND2_X1 U407 ( .A1(n468), .A2(n529), .ZN(n466) );
  NAND2_X1 U408 ( .A1(n677), .A2(n408), .ZN(n407) );
  NAND2_X1 U409 ( .A1(n347), .A2(n436), .ZN(n408) );
  NOR2_X1 U410 ( .A1(G953), .A2(G237), .ZN(n549) );
  XNOR2_X1 U411 ( .A(n428), .B(n469), .ZN(n520) );
  XNOR2_X1 U412 ( .A(G116), .B(G113), .ZN(n469) );
  XNOR2_X1 U413 ( .A(n500), .B(KEYINPUT3), .ZN(n428) );
  XNOR2_X1 U414 ( .A(G119), .B(KEYINPUT72), .ZN(n500) );
  NOR2_X1 U415 ( .A1(n690), .A2(KEYINPUT108), .ZN(n478) );
  AND2_X1 U416 ( .A1(n686), .A2(n685), .ZN(n691) );
  XNOR2_X1 U417 ( .A(n508), .B(n744), .ZN(n727) );
  XOR2_X1 U418 ( .A(KEYINPUT9), .B(G107), .Z(n560) );
  XNOR2_X1 U419 ( .A(G116), .B(G122), .ZN(n559) );
  XOR2_X1 U420 ( .A(KEYINPUT105), .B(KEYINPUT7), .Z(n563) );
  XNOR2_X1 U421 ( .A(n517), .B(n515), .ZN(n485) );
  XNOR2_X1 U422 ( .A(n514), .B(n513), .ZN(n515) );
  XNOR2_X1 U423 ( .A(n387), .B(n386), .ZN(n420) );
  NAND2_X1 U424 ( .A1(n683), .A2(n481), .ZN(n370) );
  NOR2_X1 U425 ( .A1(n575), .A2(n686), .ZN(n487) );
  INV_X1 U426 ( .A(G478), .ZN(n382) );
  OR2_X1 U427 ( .A1(n725), .A2(G902), .ZN(n383) );
  XNOR2_X1 U428 ( .A(KEYINPUT13), .B(G475), .ZN(n557) );
  NOR2_X1 U429 ( .A1(n641), .A2(n379), .ZN(n371) );
  INV_X1 U430 ( .A(G217), .ZN(n379) );
  INV_X1 U431 ( .A(n727), .ZN(n402) );
  INV_X1 U432 ( .A(G475), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n723), .B(n722), .ZN(n492) );
  INV_X1 U434 ( .A(G210), .ZN(n373) );
  NAND2_X1 U435 ( .A1(n429), .A2(n447), .ZN(n443) );
  XNOR2_X1 U436 ( .A(n523), .B(n449), .ZN(n552) );
  XNOR2_X1 U437 ( .A(KEYINPUT10), .B(G140), .ZN(n449) );
  XNOR2_X1 U438 ( .A(n415), .B(KEYINPUT65), .ZN(n521) );
  INV_X1 U439 ( .A(KEYINPUT4), .ZN(n415) );
  NAND2_X1 U440 ( .A1(n409), .A2(n410), .ZN(n404) );
  OR2_X1 U441 ( .A1(G237), .A2(G902), .ZN(n530) );
  XNOR2_X1 U442 ( .A(n746), .B(n463), .ZN(n462) );
  INV_X1 U443 ( .A(KEYINPUT76), .ZN(n463) );
  XNOR2_X1 U444 ( .A(n427), .B(G107), .ZN(n519) );
  XNOR2_X1 U445 ( .A(G104), .B(G110), .ZN(n427) );
  INV_X1 U446 ( .A(KEYINPUT95), .ZN(n513) );
  INV_X1 U447 ( .A(KEYINPUT48), .ZN(n386) );
  NOR2_X1 U448 ( .A1(n575), .A2(n480), .ZN(n476) );
  OR2_X1 U449 ( .A1(n718), .A2(G902), .ZN(n484) );
  XNOR2_X1 U450 ( .A(n533), .B(KEYINPUT19), .ZN(n534) );
  XNOR2_X1 U451 ( .A(n502), .B(n494), .ZN(n493) );
  INV_X1 U452 ( .A(KEYINPUT5), .ZN(n494) );
  INV_X1 U453 ( .A(G953), .ZN(n748) );
  XNOR2_X1 U454 ( .A(n520), .B(n424), .ZN(n736) );
  XNOR2_X1 U455 ( .A(n519), .B(n425), .ZN(n424) );
  XNOR2_X1 U456 ( .A(n426), .B(G122), .ZN(n425) );
  INV_X1 U457 ( .A(KEYINPUT16), .ZN(n426) );
  INV_X1 U458 ( .A(KEYINPUT86), .ZN(n638) );
  XNOR2_X1 U459 ( .A(n512), .B(n349), .ZN(n440) );
  XNOR2_X1 U460 ( .A(n570), .B(KEYINPUT22), .ZN(n571) );
  XNOR2_X1 U461 ( .A(n564), .B(n460), .ZN(n725) );
  XNOR2_X1 U462 ( .A(n563), .B(n562), .ZN(n564) );
  BUF_X1 U463 ( .A(G953), .Z(n381) );
  INV_X1 U464 ( .A(KEYINPUT40), .ZN(n448) );
  NAND2_X1 U465 ( .A1(n369), .A2(n368), .ZN(n367) );
  INV_X1 U466 ( .A(n614), .ZN(n368) );
  XNOR2_X1 U467 ( .A(n370), .B(n357), .ZN(n369) );
  AND2_X1 U468 ( .A1(n436), .A2(n435), .ZN(n658) );
  INV_X1 U469 ( .A(n686), .ZN(n455) );
  INV_X1 U470 ( .A(KEYINPUT122), .ZN(n399) );
  INV_X1 U471 ( .A(KEYINPUT60), .ZN(n489) );
  XNOR2_X1 U472 ( .A(n716), .B(n452), .ZN(n720) );
  XNOR2_X1 U473 ( .A(n719), .B(n717), .ZN(n452) );
  INV_X1 U474 ( .A(KEYINPUT56), .ZN(n470) );
  OR2_X1 U475 ( .A1(n455), .A2(KEYINPUT87), .ZN(n346) );
  AND2_X1 U476 ( .A1(n435), .A2(n356), .ZN(n347) );
  AND2_X1 U477 ( .A1(n455), .A2(KEYINPUT87), .ZN(n348) );
  XNOR2_X1 U478 ( .A(KEYINPUT79), .B(KEYINPUT98), .ZN(n349) );
  XOR2_X1 U479 ( .A(KEYINPUT97), .B(KEYINPUT24), .Z(n350) );
  OR2_X1 U480 ( .A1(n711), .A2(n710), .ZN(n351) );
  OR2_X1 U481 ( .A1(n610), .A2(n393), .ZN(n352) );
  AND2_X1 U482 ( .A1(n435), .A2(KEYINPUT70), .ZN(n353) );
  NAND2_X1 U483 ( .A1(n430), .A2(n346), .ZN(n354) );
  AND2_X1 U484 ( .A1(n709), .A2(n351), .ZN(n355) );
  INV_X1 U485 ( .A(KEYINPUT108), .ZN(n480) );
  AND2_X1 U486 ( .A1(KEYINPUT70), .A2(KEYINPUT47), .ZN(n356) );
  XNOR2_X1 U487 ( .A(KEYINPUT73), .B(KEYINPUT34), .ZN(n357) );
  XOR2_X1 U488 ( .A(KEYINPUT46), .B(KEYINPUT64), .Z(n358) );
  XOR2_X1 U489 ( .A(n573), .B(KEYINPUT62), .Z(n359) );
  XOR2_X1 U490 ( .A(n364), .B(n714), .Z(n360) );
  INV_X1 U491 ( .A(KEYINPUT66), .ZN(n574) );
  INV_X1 U492 ( .A(KEYINPUT47), .ZN(n410) );
  INV_X1 U493 ( .A(KEYINPUT87), .ZN(n447) );
  XOR2_X1 U494 ( .A(KEYINPUT63), .B(KEYINPUT89), .Z(n361) );
  NOR2_X1 U495 ( .A1(G952), .A2(n451), .ZN(n728) );
  INV_X1 U496 ( .A(n728), .ZN(n456) );
  INV_X1 U497 ( .A(n689), .ZN(n601) );
  INV_X1 U498 ( .A(n604), .ZN(n435) );
  XNOR2_X1 U499 ( .A(n344), .B(n574), .ZN(n362) );
  XNOR2_X1 U500 ( .A(n486), .B(KEYINPUT83), .ZN(n577) );
  XNOR2_X1 U501 ( .A(n421), .B(KEYINPUT66), .ZN(n363) );
  XNOR2_X1 U502 ( .A(n430), .B(G119), .ZN(G21) );
  XNOR2_X1 U503 ( .A(n618), .B(KEYINPUT84), .ZN(n488) );
  XNOR2_X1 U504 ( .A(n397), .B(n485), .ZN(n718) );
  XNOR2_X1 U505 ( .A(n397), .B(n493), .ZN(n573) );
  BUF_X1 U506 ( .A(n715), .Z(n364) );
  NAND2_X1 U507 ( .A1(n467), .A2(n466), .ZN(n365) );
  XNOR2_X1 U508 ( .A(n403), .B(n402), .ZN(n401) );
  NAND2_X1 U509 ( .A1(n375), .A2(n371), .ZN(n403) );
  XNOR2_X1 U510 ( .A(n482), .B(KEYINPUT120), .ZN(n712) );
  INV_X2 U511 ( .A(n707), .ZN(n641) );
  NAND2_X1 U512 ( .A1(n366), .A2(n691), .ZN(n610) );
  XNOR2_X2 U513 ( .A(n366), .B(KEYINPUT1), .ZN(n690) );
  AND2_X1 U514 ( .A1(n366), .A2(n603), .ZN(n436) );
  XNOR2_X2 U515 ( .A(n484), .B(G469), .ZN(n366) );
  NOR2_X1 U516 ( .A1(n365), .A2(n641), .ZN(n380) );
  NAND2_X1 U517 ( .A1(n375), .A2(n372), .ZN(n473) );
  NOR2_X1 U518 ( .A1(n641), .A2(n373), .ZN(n372) );
  NAND2_X1 U519 ( .A1(n375), .A2(n374), .ZN(n642) );
  NOR2_X1 U520 ( .A1(n641), .A2(n377), .ZN(n374) );
  INV_X1 U521 ( .A(n365), .ZN(n375) );
  NAND2_X1 U522 ( .A1(n375), .A2(n376), .ZN(n721) );
  NOR2_X1 U523 ( .A1(n641), .A2(n378), .ZN(n376) );
  NAND2_X1 U524 ( .A1(n380), .A2(G478), .ZN(n724) );
  NAND2_X1 U525 ( .A1(n380), .A2(G469), .ZN(n716) );
  NAND2_X1 U526 ( .A1(n401), .A2(n456), .ZN(n400) );
  NAND2_X1 U527 ( .A1(n384), .A2(n706), .ZN(n708) );
  NAND2_X1 U528 ( .A1(n729), .A2(n746), .ZN(n384) );
  XNOR2_X1 U529 ( .A(n422), .B(n417), .ZN(n416) );
  XNOR2_X1 U530 ( .A(n721), .B(n492), .ZN(n491) );
  XNOR2_X1 U531 ( .A(n414), .B(n524), .ZN(n528) );
  NAND2_X1 U532 ( .A1(n472), .A2(n456), .ZN(n471) );
  NAND2_X1 U533 ( .A1(n756), .A2(n757), .ZN(n389) );
  NAND2_X1 U534 ( .A1(n392), .A2(n613), .ZN(n623) );
  INV_X1 U535 ( .A(n673), .ZN(n391) );
  NAND2_X1 U536 ( .A1(n394), .A2(n352), .ZN(n392) );
  NAND2_X1 U537 ( .A1(n609), .A2(n612), .ZN(n393) );
  AND2_X1 U538 ( .A1(n396), .A2(n395), .ZN(n394) );
  NAND2_X1 U539 ( .A1(n611), .A2(KEYINPUT77), .ZN(n395) );
  NAND2_X1 U540 ( .A1(n610), .A2(KEYINPUT77), .ZN(n396) );
  XNOR2_X1 U541 ( .A(n398), .B(n565), .ZN(n460) );
  XNOR2_X1 U542 ( .A(n400), .B(n399), .ZN(G66) );
  NAND2_X1 U543 ( .A1(n405), .A2(n404), .ZN(n438) );
  NAND2_X1 U544 ( .A1(n407), .A2(n406), .ZN(n405) );
  NAND2_X1 U545 ( .A1(n605), .A2(KEYINPUT47), .ZN(n406) );
  NAND2_X1 U546 ( .A1(n436), .A2(n353), .ZN(n409) );
  NAND2_X1 U547 ( .A1(n411), .A2(n362), .ZN(n413) );
  XNOR2_X2 U548 ( .A(n578), .B(KEYINPUT32), .ZN(n430) );
  NAND2_X1 U549 ( .A1(n363), .A2(n348), .ZN(n412) );
  XNOR2_X1 U550 ( .A(n416), .B(n521), .ZN(n414) );
  INV_X1 U551 ( .A(n755), .ZN(n445) );
  NAND2_X1 U552 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X2 U553 ( .A(n572), .B(n571), .ZN(n576) );
  XNOR2_X1 U554 ( .A(n418), .B(n736), .ZN(n715) );
  XNOR2_X1 U555 ( .A(n528), .B(n527), .ZN(n418) );
  NAND2_X1 U556 ( .A1(n446), .A2(n445), .ZN(n434) );
  XNOR2_X1 U557 ( .A(n434), .B(n433), .ZN(n432) );
  XNOR2_X2 U558 ( .A(n419), .B(G128), .ZN(n525) );
  NAND2_X1 U559 ( .A1(n432), .A2(n594), .ZN(n431) );
  NOR2_X2 U560 ( .A1(n474), .A2(n479), .ZN(n421) );
  XNOR2_X2 U561 ( .A(KEYINPUT81), .B(KEYINPUT17), .ZN(n422) );
  INV_X1 U562 ( .A(n430), .ZN(n429) );
  NAND2_X1 U563 ( .A1(n698), .A2(n436), .ZN(n627) );
  XNOR2_X1 U564 ( .A(n437), .B(KEYINPUT75), .ZN(n622) );
  NAND2_X1 U565 ( .A1(n438), .A2(n656), .ZN(n437) );
  XNOR2_X2 U566 ( .A(n440), .B(n439), .ZN(n686) );
  NOR2_X1 U567 ( .A1(n619), .A2(n441), .ZN(n620) );
  XNOR2_X2 U568 ( .A(n465), .B(KEYINPUT88), .ZN(n441) );
  AND2_X1 U569 ( .A1(n363), .A2(n455), .ZN(n650) );
  NAND2_X1 U570 ( .A1(n354), .A2(n443), .ZN(n442) );
  XNOR2_X1 U571 ( .A(n473), .B(n360), .ZN(n472) );
  NOR2_X1 U572 ( .A1(n476), .A2(n601), .ZN(n475) );
  NAND2_X1 U573 ( .A1(n488), .A2(n487), .ZN(n486) );
  XNOR2_X1 U574 ( .A(n450), .B(n361), .ZN(G57) );
  NAND2_X1 U575 ( .A1(n457), .A2(n456), .ZN(n450) );
  BUF_X2 U576 ( .A(n748), .Z(n451) );
  XNOR2_X1 U577 ( .A(n453), .B(n507), .ZN(n508) );
  XNOR2_X1 U578 ( .A(n506), .B(n464), .ZN(n453) );
  NAND2_X1 U579 ( .A1(n462), .A2(n706), .ZN(n468) );
  XNOR2_X1 U580 ( .A(n642), .B(n359), .ZN(n457) );
  AND2_X1 U581 ( .A1(n622), .A2(n668), .ZN(n461) );
  NOR2_X2 U582 ( .A1(n589), .A2(n582), .ZN(n674) );
  NAND2_X1 U583 ( .A1(n491), .A2(n456), .ZN(n490) );
  XNOR2_X1 U584 ( .A(n490), .B(n489), .ZN(G60) );
  XNOR2_X1 U585 ( .A(n505), .B(n350), .ZN(n464) );
  NAND2_X1 U586 ( .A1(n606), .A2(n607), .ZN(n465) );
  XNOR2_X1 U587 ( .A(n532), .B(n531), .ZN(n606) );
  OR2_X2 U588 ( .A1(n705), .A2(KEYINPUT2), .ZN(n467) );
  XNOR2_X1 U589 ( .A(n471), .B(n470), .ZN(G51) );
  NAND2_X1 U590 ( .A1(n576), .A2(n575), .ZN(n592) );
  NAND2_X1 U591 ( .A1(n477), .A2(n475), .ZN(n474) );
  NAND2_X1 U592 ( .A1(n576), .A2(n478), .ZN(n477) );
  NOR2_X1 U593 ( .A1(n576), .A2(n480), .ZN(n479) );
  INV_X1 U594 ( .A(n683), .ZN(n711) );
  INV_X1 U595 ( .A(n345), .ZN(n481) );
  NAND2_X1 U596 ( .A1(n483), .A2(n355), .ZN(n482) );
  NAND2_X1 U597 ( .A1(n708), .A2(n707), .ZN(n483) );
  NAND2_X1 U598 ( .A1(n705), .A2(n640), .ZN(n707) );
  NOR2_X2 U599 ( .A1(n581), .A2(n569), .ZN(n572) );
  BUF_X1 U600 ( .A(n606), .Z(n634) );
  XNOR2_X2 U601 ( .A(n601), .B(KEYINPUT6), .ZN(n618) );
  NOR2_X1 U602 ( .A1(n671), .A2(n636), .ZN(n495) );
  AND2_X1 U603 ( .A1(n549), .A2(G214), .ZN(n496) );
  XNOR2_X1 U604 ( .A(KEYINPUT90), .B(KEYINPUT33), .ZN(n579) );
  INV_X1 U605 ( .A(n670), .ZN(n636) );
  XNOR2_X1 U606 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U607 ( .A(n550), .B(n496), .ZN(n551) );
  XNOR2_X1 U608 ( .A(n552), .B(n551), .ZN(n553) );
  INV_X1 U609 ( .A(KEYINPUT77), .ZN(n612) );
  BUF_X1 U610 ( .A(n705), .Z(n729) );
  XNOR2_X1 U611 ( .A(n519), .B(n516), .ZN(n517) );
  XOR2_X1 U612 ( .A(KEYINPUT69), .B(G101), .Z(n522) );
  XNOR2_X1 U613 ( .A(G146), .B(n522), .ZN(n499) );
  XOR2_X1 U614 ( .A(KEYINPUT71), .B(G131), .Z(n546) );
  XOR2_X1 U615 ( .A(n521), .B(G137), .Z(n498) );
  NAND2_X1 U616 ( .A1(n549), .A2(G210), .ZN(n501) );
  XNOR2_X1 U617 ( .A(n520), .B(n501), .ZN(n502) );
  XOR2_X1 U618 ( .A(G137), .B(G128), .Z(n504) );
  XNOR2_X1 U619 ( .A(G119), .B(G110), .ZN(n503) );
  XNOR2_X1 U620 ( .A(n504), .B(n503), .ZN(n506) );
  XOR2_X1 U621 ( .A(KEYINPUT23), .B(KEYINPUT96), .Z(n505) );
  NAND2_X1 U622 ( .A1(G221), .A2(n561), .ZN(n507) );
  INV_X1 U623 ( .A(n552), .ZN(n744) );
  XOR2_X1 U624 ( .A(KEYINPUT25), .B(KEYINPUT99), .Z(n511) );
  INV_X1 U625 ( .A(n529), .ZN(n637) );
  NAND2_X1 U626 ( .A1(G234), .A2(n637), .ZN(n509) );
  XNOR2_X1 U627 ( .A(KEYINPUT20), .B(n509), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n566), .A2(G217), .ZN(n510) );
  XNOR2_X1 U629 ( .A(n511), .B(n510), .ZN(n512) );
  NAND2_X1 U630 ( .A1(G227), .A2(n451), .ZN(n514) );
  XNOR2_X1 U631 ( .A(G140), .B(KEYINPUT80), .ZN(n516) );
  NAND2_X1 U632 ( .A1(n530), .A2(G214), .ZN(n518) );
  XOR2_X1 U633 ( .A(KEYINPUT91), .B(n518), .Z(n607) );
  XNOR2_X1 U634 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U635 ( .A(n525), .B(KEYINPUT82), .ZN(n526) );
  XNOR2_X1 U636 ( .A(n526), .B(KEYINPUT18), .ZN(n527) );
  NOR2_X1 U637 ( .A1(n715), .A2(n529), .ZN(n532) );
  NAND2_X1 U638 ( .A1(G210), .A2(n530), .ZN(n531) );
  XOR2_X1 U639 ( .A(KEYINPUT78), .B(KEYINPUT68), .Z(n533) );
  NAND2_X1 U640 ( .A1(G234), .A2(G237), .ZN(n535) );
  XNOR2_X1 U641 ( .A(n535), .B(KEYINPUT14), .ZN(n538) );
  NAND2_X1 U642 ( .A1(n538), .A2(G952), .ZN(n536) );
  XOR2_X1 U643 ( .A(KEYINPUT92), .B(n536), .Z(n703) );
  NAND2_X1 U644 ( .A1(n451), .A2(n703), .ZN(n599) );
  INV_X1 U645 ( .A(n599), .ZN(n541) );
  NOR2_X1 U646 ( .A1(G898), .A2(n451), .ZN(n537) );
  XNOR2_X1 U647 ( .A(KEYINPUT93), .B(n537), .ZN(n740) );
  NAND2_X1 U648 ( .A1(G902), .A2(n538), .ZN(n596) );
  NOR2_X1 U649 ( .A1(n740), .A2(n596), .ZN(n539) );
  XNOR2_X1 U650 ( .A(n539), .B(KEYINPUT94), .ZN(n540) );
  NOR2_X1 U651 ( .A1(n541), .A2(n540), .ZN(n542) );
  INV_X1 U652 ( .A(KEYINPUT0), .ZN(n543) );
  XNOR2_X1 U653 ( .A(n545), .B(n544), .ZN(n556) );
  XNOR2_X1 U654 ( .A(n546), .B(KEYINPUT102), .ZN(n554) );
  XOR2_X1 U655 ( .A(KEYINPUT104), .B(KEYINPUT12), .Z(n548) );
  XNOR2_X1 U656 ( .A(KEYINPUT103), .B(KEYINPUT11), .ZN(n547) );
  XNOR2_X1 U657 ( .A(n548), .B(n547), .ZN(n550) );
  XNOR2_X1 U658 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U659 ( .A(n556), .B(n555), .ZN(n723) );
  NOR2_X1 U660 ( .A1(G902), .A2(n723), .ZN(n558) );
  XNOR2_X1 U661 ( .A(n560), .B(n559), .ZN(n565) );
  NAND2_X1 U662 ( .A1(G217), .A2(n561), .ZN(n562) );
  INV_X1 U663 ( .A(n588), .ZN(n582) );
  NAND2_X1 U664 ( .A1(n566), .A2(G221), .ZN(n567) );
  XOR2_X1 U665 ( .A(KEYINPUT21), .B(n567), .Z(n685) );
  NAND2_X1 U666 ( .A1(n674), .A2(n685), .ZN(n568) );
  XOR2_X1 U667 ( .A(KEYINPUT107), .B(n568), .Z(n569) );
  XOR2_X1 U668 ( .A(KEYINPUT67), .B(KEYINPUT74), .Z(n570) );
  NAND2_X1 U669 ( .A1(n690), .A2(n691), .ZN(n584) );
  OR2_X1 U670 ( .A1(n618), .A2(n584), .ZN(n580) );
  NAND2_X1 U671 ( .A1(n589), .A2(n582), .ZN(n614) );
  NOR2_X1 U672 ( .A1(n345), .A2(n610), .ZN(n583) );
  NAND2_X1 U673 ( .A1(n689), .A2(n583), .ZN(n646) );
  NOR2_X1 U674 ( .A1(n689), .A2(n584), .ZN(n696) );
  NAND2_X1 U675 ( .A1(n481), .A2(n696), .ZN(n585) );
  XNOR2_X1 U676 ( .A(n585), .B(KEYINPUT101), .ZN(n586) );
  XNOR2_X1 U677 ( .A(KEYINPUT31), .B(n586), .ZN(n663) );
  NAND2_X1 U678 ( .A1(n646), .A2(n663), .ZN(n590) );
  NOR2_X1 U679 ( .A1(n589), .A2(n588), .ZN(n587) );
  XOR2_X1 U680 ( .A(KEYINPUT106), .B(n587), .Z(n664) );
  NAND2_X1 U681 ( .A1(n589), .A2(n588), .ZN(n624) );
  NAND2_X1 U682 ( .A1(n664), .A2(n624), .ZN(n677) );
  AND2_X1 U683 ( .A1(n590), .A2(n677), .ZN(n593) );
  NAND2_X1 U684 ( .A1(n686), .A2(n618), .ZN(n591) );
  NOR2_X1 U685 ( .A1(n592), .A2(n591), .ZN(n643) );
  NOR2_X1 U686 ( .A1(n593), .A2(n643), .ZN(n594) );
  INV_X1 U687 ( .A(n677), .ZN(n605) );
  NOR2_X1 U688 ( .A1(G900), .A2(n596), .ZN(n597) );
  NAND2_X1 U689 ( .A1(n381), .A2(n597), .ZN(n598) );
  NAND2_X1 U690 ( .A1(n599), .A2(n598), .ZN(n609) );
  NAND2_X1 U691 ( .A1(n685), .A2(n609), .ZN(n600) );
  NOR2_X1 U692 ( .A1(n686), .A2(n600), .ZN(n616) );
  AND2_X1 U693 ( .A1(n601), .A2(n616), .ZN(n602) );
  XNOR2_X1 U694 ( .A(KEYINPUT28), .B(n602), .ZN(n603) );
  INV_X1 U695 ( .A(n607), .ZN(n672) );
  NOR2_X1 U696 ( .A1(n672), .A2(n689), .ZN(n608) );
  XNOR2_X1 U697 ( .A(KEYINPUT30), .B(n608), .ZN(n613) );
  INV_X1 U698 ( .A(n609), .ZN(n611) );
  NOR2_X1 U699 ( .A1(n614), .A2(n623), .ZN(n615) );
  NAND2_X1 U700 ( .A1(n634), .A2(n615), .ZN(n656) );
  XNOR2_X1 U701 ( .A(KEYINPUT109), .B(n624), .ZN(n657) );
  NAND2_X1 U702 ( .A1(n616), .A2(n657), .ZN(n617) );
  NOR2_X1 U703 ( .A1(n618), .A2(n617), .ZN(n630) );
  INV_X1 U704 ( .A(n630), .ZN(n619) );
  XNOR2_X1 U705 ( .A(KEYINPUT36), .B(n620), .ZN(n621) );
  NAND2_X1 U706 ( .A1(n621), .A2(n690), .ZN(n668) );
  XNOR2_X1 U707 ( .A(KEYINPUT38), .B(n634), .ZN(n673) );
  XOR2_X1 U708 ( .A(KEYINPUT111), .B(KEYINPUT42), .Z(n628) );
  NOR2_X1 U709 ( .A1(n672), .A2(n673), .ZN(n678) );
  NAND2_X1 U710 ( .A1(n674), .A2(n678), .ZN(n626) );
  XNOR2_X1 U711 ( .A(KEYINPUT41), .B(n626), .ZN(n698) );
  INV_X1 U712 ( .A(n698), .ZN(n710) );
  XNOR2_X1 U713 ( .A(n628), .B(n627), .ZN(n757) );
  NOR2_X1 U714 ( .A1(n690), .A2(n672), .ZN(n629) );
  NAND2_X1 U715 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U716 ( .A(KEYINPUT110), .B(n631), .ZN(n632) );
  XOR2_X1 U717 ( .A(KEYINPUT43), .B(n632), .Z(n633) );
  NOR2_X1 U718 ( .A1(n634), .A2(n633), .ZN(n671) );
  OR2_X1 U719 ( .A1(n635), .A2(n664), .ZN(n670) );
  INV_X1 U720 ( .A(KEYINPUT2), .ZN(n706) );
  NAND2_X1 U721 ( .A1(n746), .A2(KEYINPUT2), .ZN(n639) );
  XOR2_X1 U722 ( .A(G101), .B(n643), .Z(G3) );
  INV_X1 U723 ( .A(n657), .ZN(n661) );
  NOR2_X1 U724 ( .A1(n646), .A2(n661), .ZN(n644) );
  XOR2_X1 U725 ( .A(KEYINPUT112), .B(n644), .Z(n645) );
  XNOR2_X1 U726 ( .A(G104), .B(n645), .ZN(G6) );
  NOR2_X1 U727 ( .A1(n664), .A2(n646), .ZN(n648) );
  XNOR2_X1 U728 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n647) );
  XNOR2_X1 U729 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U730 ( .A(G107), .B(n649), .ZN(G9) );
  XOR2_X1 U731 ( .A(n650), .B(G110), .Z(G12) );
  XOR2_X1 U732 ( .A(KEYINPUT114), .B(KEYINPUT29), .Z(n653) );
  INV_X1 U733 ( .A(n664), .ZN(n651) );
  NAND2_X1 U734 ( .A1(n658), .A2(n651), .ZN(n652) );
  XNOR2_X1 U735 ( .A(n653), .B(n652), .ZN(n655) );
  XOR2_X1 U736 ( .A(G128), .B(KEYINPUT113), .Z(n654) );
  XNOR2_X1 U737 ( .A(n655), .B(n654), .ZN(G30) );
  XNOR2_X1 U738 ( .A(G143), .B(n656), .ZN(G45) );
  XOR2_X1 U739 ( .A(G146), .B(KEYINPUT115), .Z(n660) );
  NAND2_X1 U740 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U741 ( .A(n660), .B(n659), .ZN(G48) );
  NOR2_X1 U742 ( .A1(n663), .A2(n661), .ZN(n662) );
  XOR2_X1 U743 ( .A(G113), .B(n662), .Z(G15) );
  NOR2_X1 U744 ( .A1(n664), .A2(n663), .ZN(n665) );
  XOR2_X1 U745 ( .A(KEYINPUT116), .B(n665), .Z(n666) );
  XNOR2_X1 U746 ( .A(G116), .B(n666), .ZN(G18) );
  XOR2_X1 U747 ( .A(G125), .B(KEYINPUT37), .Z(n667) );
  XNOR2_X1 U748 ( .A(n668), .B(n667), .ZN(G27) );
  XOR2_X1 U749 ( .A(G134), .B(KEYINPUT117), .Z(n669) );
  XNOR2_X1 U750 ( .A(n670), .B(n669), .ZN(G36) );
  XOR2_X1 U751 ( .A(G140), .B(n671), .Z(G42) );
  AND2_X1 U752 ( .A1(n673), .A2(n672), .ZN(n676) );
  INV_X1 U753 ( .A(n674), .ZN(n675) );
  NOR2_X1 U754 ( .A1(n676), .A2(n675), .ZN(n681) );
  NAND2_X1 U755 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U756 ( .A(KEYINPUT118), .B(n679), .Z(n680) );
  NOR2_X1 U757 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U758 ( .A(n682), .B(KEYINPUT119), .ZN(n684) );
  NAND2_X1 U759 ( .A1(n684), .A2(n683), .ZN(n701) );
  NOR2_X1 U760 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U761 ( .A(n687), .B(KEYINPUT49), .ZN(n688) );
  NAND2_X1 U762 ( .A1(n689), .A2(n688), .ZN(n694) );
  NOR2_X1 U763 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U764 ( .A(n692), .B(KEYINPUT50), .ZN(n693) );
  NOR2_X1 U765 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U766 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U767 ( .A(KEYINPUT51), .B(n697), .ZN(n699) );
  NAND2_X1 U768 ( .A1(n699), .A2(n698), .ZN(n700) );
  NAND2_X1 U769 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U770 ( .A(n702), .B(KEYINPUT52), .ZN(n704) );
  NAND2_X1 U771 ( .A1(n704), .A2(n703), .ZN(n709) );
  XNOR2_X1 U772 ( .A(n713), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U773 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n714) );
  XOR2_X1 U774 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n717) );
  BUF_X1 U775 ( .A(n718), .Z(n719) );
  NOR2_X1 U776 ( .A1(n728), .A2(n720), .ZN(G54) );
  XOR2_X1 U777 ( .A(KEYINPUT59), .B(KEYINPUT121), .Z(n722) );
  XNOR2_X1 U778 ( .A(n725), .B(n724), .ZN(n726) );
  NOR2_X1 U779 ( .A1(n728), .A2(n726), .ZN(G63) );
  NAND2_X1 U780 ( .A1(n729), .A2(n451), .ZN(n730) );
  XNOR2_X1 U781 ( .A(n730), .B(KEYINPUT124), .ZN(n735) );
  XOR2_X1 U782 ( .A(KEYINPUT61), .B(KEYINPUT123), .Z(n732) );
  NAND2_X1 U783 ( .A1(G224), .A2(n381), .ZN(n731) );
  XNOR2_X1 U784 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U785 ( .A1(n733), .A2(G898), .ZN(n734) );
  NAND2_X1 U786 ( .A1(n735), .A2(n734), .ZN(n742) );
  XOR2_X1 U787 ( .A(KEYINPUT126), .B(KEYINPUT125), .Z(n738) );
  XNOR2_X1 U788 ( .A(n736), .B(G101), .ZN(n737) );
  XNOR2_X1 U789 ( .A(n738), .B(n737), .ZN(n739) );
  NAND2_X1 U790 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U791 ( .A(n742), .B(n741), .Z(G69) );
  XNOR2_X1 U792 ( .A(n743), .B(KEYINPUT127), .ZN(n745) );
  XOR2_X1 U793 ( .A(n745), .B(n744), .Z(n750) );
  INV_X1 U794 ( .A(n750), .ZN(n747) );
  XNOR2_X1 U795 ( .A(n747), .B(n746), .ZN(n749) );
  NAND2_X1 U796 ( .A1(n749), .A2(n451), .ZN(n754) );
  XNOR2_X1 U797 ( .A(G227), .B(n750), .ZN(n751) );
  NAND2_X1 U798 ( .A1(n751), .A2(G900), .ZN(n752) );
  NAND2_X1 U799 ( .A1(n752), .A2(n381), .ZN(n753) );
  NAND2_X1 U800 ( .A1(n754), .A2(n753), .ZN(G72) );
  XOR2_X1 U801 ( .A(n755), .B(G122), .Z(G24) );
  XNOR2_X1 U802 ( .A(n756), .B(G131), .ZN(G33) );
  XNOR2_X1 U803 ( .A(G137), .B(n757), .ZN(G39) );
endmodule

