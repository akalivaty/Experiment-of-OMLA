//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 1 1 0 0 1 0 1 1 0 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  AND2_X1   g001(.A1(KEYINPUT64), .A2(G143), .ZN(new_n188));
  NOR2_X1   g002(.A1(KEYINPUT64), .A2(G143), .ZN(new_n189));
  OAI21_X1  g003(.A(G146), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G146), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G128), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n194), .A2(KEYINPUT1), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n190), .A2(new_n193), .A3(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT67), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT67), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n190), .A2(new_n198), .A3(new_n193), .A4(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  NOR3_X1   g014(.A1(new_n188), .A2(new_n189), .A3(G146), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT1), .ZN(new_n202));
  OAI21_X1  g016(.A(G128), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n190), .A2(new_n193), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n200), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT84), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G107), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n208), .A2(G107), .ZN(new_n210));
  INV_X1    g024(.A(G107), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT84), .A3(G104), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n210), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G101), .ZN(new_n214));
  OAI21_X1  g028(.A(KEYINPUT3), .B1(new_n208), .B2(G107), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT3), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n216), .A2(new_n211), .A3(G104), .ZN(new_n217));
  INV_X1    g031(.A(G101), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n215), .A2(new_n217), .A3(new_n218), .A4(new_n210), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n206), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(G128), .B1(new_n192), .B2(new_n202), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT65), .B1(new_n224), .B2(G143), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n191), .A3(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n223), .B1(new_n201), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT68), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n231), .B(new_n223), .C1(new_n201), .C2(new_n228), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n200), .A2(new_n230), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n220), .A2(KEYINPUT85), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT85), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n214), .A2(new_n235), .A3(new_n219), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n222), .B1(new_n233), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n239));
  INV_X1    g053(.A(G137), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(G134), .ZN(new_n241));
  INV_X1    g055(.A(G134), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT66), .A3(G137), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT11), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n245), .B1(new_n242), .B2(G137), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n242), .A2(G137), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT11), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n244), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G131), .ZN(new_n250));
  INV_X1    g064(.A(G131), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n244), .A2(new_n248), .A3(new_n251), .A4(new_n246), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n238), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT12), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n233), .A2(new_n237), .A3(KEYINPUT10), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT86), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT10), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n257), .A2(new_n258), .B1(new_n222), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n253), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n219), .A2(KEYINPUT4), .ZN(new_n262));
  NAND3_X1  g076(.A1(new_n215), .A2(new_n217), .A3(new_n210), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G101), .ZN(new_n264));
  XNOR2_X1  g078(.A(new_n262), .B(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n266));
  XOR2_X1   g080(.A(KEYINPUT0), .B(G128), .Z(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n201), .B2(new_n228), .ZN(new_n268));
  NAND4_X1  g082(.A1(new_n190), .A2(KEYINPUT0), .A3(G128), .A4(new_n193), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n266), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND3_X1   g084(.A1(new_n268), .A2(new_n266), .A3(new_n269), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n265), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n233), .A2(new_n237), .A3(KEYINPUT86), .A4(KEYINPUT10), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n260), .A2(new_n261), .A3(new_n272), .A4(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n256), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(G110), .B(G140), .ZN(new_n276));
  INV_X1    g090(.A(G227), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(G953), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n276), .B(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n274), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n281), .A2(new_n279), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n200), .A2(new_n230), .A3(new_n232), .ZN(new_n283));
  INV_X1    g097(.A(new_n236), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n235), .B1(new_n214), .B2(new_n219), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT10), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n258), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n222), .A2(new_n259), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n287), .A2(new_n288), .A3(new_n272), .A4(new_n273), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(new_n253), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n282), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n280), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n187), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n290), .A2(new_n274), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n279), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(KEYINPUT88), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n282), .A2(new_n256), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT88), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n295), .A2(new_n299), .A3(new_n279), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n297), .A2(new_n298), .A3(new_n300), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT87), .B(G469), .Z(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n293), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT89), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n301), .A2(KEYINPUT89), .A3(new_n293), .A4(new_n302), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n294), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G221), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT9), .B(G234), .Z(new_n309));
  AOI21_X1  g123(.A(new_n308), .B1(new_n309), .B2(new_n293), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g125(.A(G214), .B1(G237), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g127(.A1(KEYINPUT2), .A2(G113), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT70), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT70), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n316), .B1(KEYINPUT2), .B2(G113), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(KEYINPUT2), .A2(G113), .ZN(new_n319));
  XNOR2_X1  g133(.A(G116), .B(G119), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT5), .ZN(new_n322));
  INV_X1    g136(.A(G119), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(G116), .ZN(new_n324));
  XNOR2_X1  g138(.A(new_n324), .B(KEYINPUT90), .ZN(new_n325));
  INV_X1    g139(.A(new_n320), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n325), .B(G113), .C1(new_n322), .C2(new_n326), .ZN(new_n327));
  AND3_X1   g141(.A1(new_n237), .A2(new_n321), .A3(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT91), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n318), .A2(new_n319), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n326), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n321), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n265), .A2(new_n333), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n327), .A2(new_n321), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n237), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT91), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n330), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  XOR2_X1   g152(.A(G110), .B(G122), .Z(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n339), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n330), .A2(new_n341), .A3(new_n337), .A4(new_n334), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(KEYINPUT6), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT6), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n338), .A2(new_n344), .A3(new_n339), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n268), .A2(new_n269), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G125), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n347), .B1(new_n233), .B2(G125), .ZN(new_n348));
  INV_X1    g162(.A(G953), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G224), .ZN(new_n350));
  XOR2_X1   g164(.A(new_n348), .B(new_n350), .Z(new_n351));
  NAND3_X1  g165(.A1(new_n343), .A2(new_n345), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(KEYINPUT7), .ZN(new_n353));
  XOR2_X1   g167(.A(new_n348), .B(new_n353), .Z(new_n354));
  XOR2_X1   g168(.A(new_n339), .B(KEYINPUT8), .Z(new_n355));
  NOR2_X1   g169(.A1(new_n335), .A2(new_n221), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n355), .B1(new_n328), .B2(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n354), .A2(new_n342), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n352), .A2(new_n293), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(G210), .B1(G237), .B2(G902), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n361), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n313), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G237), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n191), .A2(new_n365), .A3(new_n349), .A4(G214), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT64), .B(G143), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n365), .A2(new_n349), .A3(G214), .ZN(new_n368));
  OAI211_X1 g182(.A(G131), .B(new_n366), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(KEYINPUT93), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT17), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(new_n251), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT95), .ZN(new_n375));
  OR2_X1    g189(.A1(new_n370), .A2(new_n371), .ZN(new_n376));
  XNOR2_X1  g190(.A(G125), .B(G140), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(KEYINPUT16), .ZN(new_n378));
  INV_X1    g192(.A(G125), .ZN(new_n379));
  OR3_X1    g193(.A1(new_n379), .A2(KEYINPUT16), .A3(G140), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(G146), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT95), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n370), .A2(new_n383), .A3(new_n371), .A4(new_n373), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n375), .A2(new_n376), .A3(new_n382), .A4(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT18), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n372), .B1(new_n386), .B2(new_n251), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n377), .B(new_n224), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n387), .B(new_n388), .C1(new_n386), .C2(new_n369), .ZN(new_n389));
  XNOR2_X1  g203(.A(G113), .B(G122), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(new_n208), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(KEYINPUT94), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n385), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n370), .A2(new_n373), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n378), .A2(G146), .A3(new_n380), .ZN(new_n396));
  XOR2_X1   g210(.A(new_n377), .B(KEYINPUT19), .Z(new_n397));
  OAI21_X1  g211(.A(new_n396), .B1(new_n397), .B2(G146), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n389), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n391), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(G475), .B1(new_n394), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n293), .ZN(new_n403));
  XNOR2_X1  g217(.A(KEYINPUT92), .B(KEYINPUT20), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n405), .B1(KEYINPUT20), .B2(new_n403), .ZN(new_n406));
  INV_X1    g220(.A(new_n394), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n391), .B1(new_n385), .B2(new_n389), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n293), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(KEYINPUT96), .B(G475), .Z(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n406), .A2(new_n411), .ZN(new_n412));
  XOR2_X1   g226(.A(KEYINPUT21), .B(G898), .Z(new_n413));
  XNOR2_X1  g227(.A(new_n413), .B(KEYINPUT98), .ZN(new_n414));
  AOI211_X1 g228(.A(new_n293), .B(new_n349), .C1(G234), .C2(G237), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G952), .ZN(new_n417));
  AOI211_X1 g231(.A(G953), .B(new_n417), .C1(G234), .C2(G237), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(KEYINPUT99), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT97), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT15), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G478), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n309), .A2(G217), .A3(new_n349), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n367), .A2(G128), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n428), .B1(G128), .B2(new_n191), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(G134), .ZN(new_n430));
  INV_X1    g244(.A(G116), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(KEYINPUT14), .A3(G122), .ZN(new_n432));
  XNOR2_X1  g246(.A(G116), .B(G122), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(G107), .B(new_n432), .C1(new_n434), .C2(KEYINPUT14), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n430), .B(new_n435), .C1(G107), .C2(new_n434), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT13), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n367), .A2(new_n437), .A3(G128), .ZN(new_n438));
  OAI211_X1 g252(.A(G134), .B(new_n438), .C1(new_n429), .C2(new_n437), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n433), .B(new_n211), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n439), .B(new_n440), .C1(G134), .C2(new_n429), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n427), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n436), .A2(new_n441), .A3(new_n427), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n425), .B1(new_n445), .B2(new_n293), .ZN(new_n446));
  INV_X1    g260(.A(new_n444), .ZN(new_n447));
  OAI211_X1 g261(.A(new_n293), .B(new_n425), .C1(new_n447), .C2(new_n442), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n423), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n447), .A2(new_n442), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n424), .B(G478), .C1(new_n451), .C2(G902), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(KEYINPUT97), .A3(new_n448), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n412), .A2(new_n422), .A3(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n311), .A2(new_n364), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT100), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n323), .A2(G128), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n194), .A2(G119), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  XOR2_X1   g275(.A(KEYINPUT24), .B(G110), .Z(new_n462));
  AOI21_X1  g276(.A(new_n382), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT23), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n459), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n194), .A2(KEYINPUT23), .A3(G119), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n465), .A2(new_n458), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G110), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  XOR2_X1   g283(.A(KEYINPUT81), .B(G110), .Z(new_n470));
  OAI22_X1  g284(.A1(new_n467), .A2(new_n470), .B1(new_n461), .B2(new_n462), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n377), .A2(new_n224), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n471), .A2(new_n396), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g288(.A(KEYINPUT22), .B(G137), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n349), .A2(G221), .A3(G234), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n475), .B(new_n476), .Z(new_n477));
  XNOR2_X1  g291(.A(new_n474), .B(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT82), .B1(new_n479), .B2(G902), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n480), .B(KEYINPUT25), .ZN(new_n481));
  INV_X1    g295(.A(G217), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(G234), .B2(new_n293), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n483), .A2(G902), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n485), .B(KEYINPUT83), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n478), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n240), .A2(G134), .ZN(new_n489));
  OAI21_X1  g303(.A(G131), .B1(new_n247), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n252), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n233), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT69), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT30), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n261), .A2(new_n346), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT69), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n233), .A2(new_n498), .A3(new_n492), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n494), .A2(new_n495), .A3(new_n497), .A4(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n253), .B1(new_n271), .B2(new_n270), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT72), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n253), .B(KEYINPUT72), .C1(new_n271), .C2(new_n270), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT73), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n491), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n252), .A2(KEYINPUT73), .A3(new_n490), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g322(.A1(new_n503), .A2(new_n504), .B1(new_n233), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n500), .B1(new_n509), .B2(new_n495), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n333), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT31), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n503), .A2(new_n504), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT74), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n320), .B1(new_n318), .B2(new_n319), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n332), .A2(KEYINPUT74), .A3(new_n321), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n508), .B2(new_n233), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n513), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT75), .B(KEYINPUT27), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n365), .A2(new_n349), .A3(G210), .ZN(new_n523));
  XNOR2_X1  g337(.A(new_n522), .B(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(KEYINPUT26), .B(G101), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n524), .B(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n511), .A2(new_n512), .A3(new_n521), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(KEYINPUT76), .ZN(new_n529));
  AND2_X1   g343(.A1(new_n513), .A2(new_n520), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n530), .B1(new_n510), .B2(new_n333), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT76), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n512), .A4(new_n527), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n233), .A2(new_n498), .A3(new_n492), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n498), .B1(new_n233), .B2(new_n492), .ZN(new_n536));
  NOR3_X1   g350(.A1(new_n535), .A2(new_n536), .A3(new_n496), .ZN(new_n537));
  INV_X1    g351(.A(new_n333), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n521), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT28), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n508), .A2(new_n233), .ZN(new_n541));
  INV_X1    g355(.A(new_n519), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n501), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT77), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT28), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n544), .B1(new_n543), .B2(new_n545), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n527), .B1(new_n540), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n511), .A2(new_n521), .A3(new_n527), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n549), .A2(KEYINPUT78), .B1(new_n550), .B2(KEYINPUT31), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n494), .A2(new_n497), .A3(new_n499), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n333), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n545), .B1(new_n553), .B2(new_n521), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n543), .A2(new_n545), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT77), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n526), .B1(new_n554), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT78), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n534), .A2(new_n551), .A3(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(G472), .A2(G902), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n562), .A2(KEYINPUT32), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT80), .ZN(new_n565));
  INV_X1    g379(.A(new_n563), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n550), .A2(KEYINPUT31), .ZN(new_n567));
  OAI211_X1 g381(.A(KEYINPUT78), .B(new_n526), .C1(new_n554), .C2(new_n558), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n561), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n566), .B1(new_n569), .B2(new_n534), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT80), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n571), .A3(KEYINPUT32), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n565), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n562), .A2(new_n563), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT32), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n531), .A2(new_n526), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n527), .B1(new_n554), .B2(new_n558), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT29), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n542), .B1(new_n513), .B2(new_n541), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT28), .B1(new_n530), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT79), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n581), .B1(new_n546), .B2(new_n547), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n556), .A2(KEYINPUT79), .A3(new_n557), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT29), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n526), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n293), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  OR2_X1    g402(.A1(new_n578), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g403(.A1(new_n574), .A2(new_n575), .B1(G472), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n488), .B1(new_n573), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n359), .B(new_n361), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n312), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n307), .A2(new_n593), .A3(new_n310), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT100), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n594), .A2(new_n595), .A3(new_n455), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n457), .A2(new_n591), .A3(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(KEYINPUT101), .B(G101), .Z(new_n598));
  XNOR2_X1  g412(.A(new_n597), .B(new_n598), .ZN(G3));
  OR2_X1    g413(.A1(new_n307), .A2(new_n310), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n600), .A2(new_n488), .ZN(new_n601));
  INV_X1    g415(.A(new_n412), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n451), .A2(G902), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(G478), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n451), .B1(KEYINPUT102), .B2(KEYINPUT33), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n605), .B1(KEYINPUT102), .B2(KEYINPUT33), .ZN(new_n606));
  OR3_X1    g420(.A1(new_n445), .A2(KEYINPUT102), .A3(KEYINPUT33), .ZN(new_n607));
  AOI21_X1  g421(.A(G902), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n604), .B1(new_n608), .B2(G478), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n364), .A2(new_n421), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n562), .A2(new_n293), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(G472), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n616), .A2(new_n570), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n601), .A2(new_n613), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G104), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT103), .B(KEYINPUT34), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G6));
  INV_X1    g435(.A(KEYINPUT104), .ZN(new_n622));
  INV_X1    g436(.A(new_n404), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n402), .A2(new_n293), .A3(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n405), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n625), .A2(new_n454), .A3(new_n411), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n622), .B1(new_n626), .B2(new_n422), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n405), .A2(new_n624), .B1(new_n409), .B2(new_n410), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n628), .A2(KEYINPUT104), .A3(new_n421), .A4(new_n454), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n627), .A2(new_n364), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(KEYINPUT105), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT105), .ZN(new_n632));
  NAND4_X1  g446(.A1(new_n627), .A2(new_n364), .A3(new_n632), .A4(new_n629), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n601), .A2(new_n634), .A3(new_n617), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT35), .B(G107), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G9));
  INV_X1    g451(.A(new_n477), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n638), .A2(KEYINPUT36), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n474), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n486), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n484), .A2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n457), .A2(new_n596), .A3(new_n617), .A4(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  AOI21_X1  g459(.A(new_n571), .B1(new_n570), .B2(KEYINPUT32), .ZN(new_n646));
  AND4_X1   g460(.A1(new_n571), .A2(new_n562), .A3(KEYINPUT32), .A4(new_n563), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n590), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n418), .B1(new_n415), .B2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n626), .A2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n648), .A2(new_n594), .A3(new_n642), .A4(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT106), .ZN(new_n653));
  INV_X1    g467(.A(new_n642), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n573), .B2(new_n590), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n655), .A2(new_n656), .A3(new_n594), .A4(new_n651), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n653), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(G128), .ZN(G30));
  NAND2_X1  g473(.A1(new_n574), .A2(new_n575), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n531), .A2(new_n526), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n521), .B1(new_n509), .B2(new_n542), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n293), .B1(new_n662), .B2(new_n527), .ZN(new_n663));
  OAI21_X1  g477(.A(G472), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n573), .A2(new_n660), .A3(new_n664), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n412), .A2(new_n312), .A3(new_n454), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n592), .B(KEYINPUT38), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n665), .A2(new_n654), .A3(new_n666), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT107), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n650), .B(KEYINPUT39), .Z(new_n670));
  NAND2_X1  g484(.A1(new_n311), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n671), .B(KEYINPUT40), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(new_n367), .Z(G45));
  INV_X1    g488(.A(new_n650), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n610), .A2(new_n675), .ZN(new_n676));
  INV_X1    g490(.A(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n655), .A2(new_n594), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  NAND2_X1  g493(.A1(new_n305), .A2(new_n306), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n301), .A2(new_n293), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(G469), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n310), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n591), .A2(new_n613), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  NAND3_X1  g501(.A1(new_n591), .A2(new_n634), .A3(new_n684), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G116), .ZN(G18));
  NOR3_X1   g503(.A1(new_n683), .A2(new_n593), .A3(new_n310), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n655), .A2(new_n455), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G119), .ZN(G21));
  AND2_X1   g506(.A1(new_n666), .A2(new_n592), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n693), .A2(new_n421), .ZN(new_n694));
  INV_X1    g508(.A(new_n488), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n526), .A2(new_n584), .B1(new_n550), .B2(KEYINPUT31), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n534), .B1(new_n696), .B2(KEYINPUT108), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n584), .A2(new_n526), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n567), .A3(KEYINPUT108), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n563), .B1(new_n697), .B2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n698), .A2(new_n567), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(new_n534), .A3(new_n699), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(KEYINPUT109), .A3(new_n563), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n616), .B1(new_n703), .B2(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n694), .A2(new_n695), .A3(new_n709), .A4(new_n684), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  AOI22_X1  g525(.A1(new_n704), .A2(new_n705), .B1(new_n533), .B2(new_n529), .ZN(new_n712));
  AOI211_X1 g526(.A(new_n702), .B(new_n566), .C1(new_n712), .C2(new_n699), .ZN(new_n713));
  AOI21_X1  g527(.A(KEYINPUT109), .B1(new_n707), .B2(new_n563), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n615), .B(new_n642), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT110), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n703), .A2(new_n708), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT110), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n717), .A2(new_n718), .A3(new_n615), .A4(new_n642), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n720), .A2(new_n677), .A3(new_n690), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  INV_X1    g536(.A(new_n590), .ZN(new_n723));
  INV_X1    g537(.A(new_n564), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n695), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n592), .A2(new_n313), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n311), .A2(new_n610), .A3(new_n675), .A4(new_n726), .ZN(new_n727));
  OAI21_X1  g541(.A(KEYINPUT42), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n676), .A2(KEYINPUT42), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n591), .A2(new_n311), .A3(new_n726), .A4(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n728), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n251), .ZN(G33));
  NAND4_X1  g546(.A1(new_n591), .A2(new_n311), .A3(new_n651), .A4(new_n726), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G134), .ZN(G36));
  INV_X1    g548(.A(KEYINPUT45), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n292), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n280), .A2(KEYINPUT45), .A3(new_n291), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n736), .A2(G469), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(G469), .A2(G902), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT46), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n740), .B(KEYINPUT111), .Z(new_n741));
  NAND3_X1  g555(.A1(new_n738), .A2(KEYINPUT46), .A3(new_n739), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n742), .A2(new_n680), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n310), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n670), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT44), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n617), .A2(new_n654), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT115), .ZN(new_n750));
  INV_X1    g564(.A(new_n609), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(KEYINPUT43), .A3(new_n602), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT114), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n751), .A2(KEYINPUT113), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n751), .A2(KEYINPUT113), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n755), .A2(new_n602), .A3(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n754), .B1(new_n757), .B2(KEYINPUT43), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n750), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n747), .B1(new_n748), .B2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n748), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n726), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(new_n240), .ZN(G39));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n744), .B(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n573), .A2(new_n590), .A3(new_n488), .A4(new_n726), .ZN(new_n767));
  OR3_X1    g581(.A1(new_n766), .A2(new_n676), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  AND2_X1   g583(.A1(new_n709), .A2(new_n695), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n758), .A2(new_n418), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n683), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n310), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n771), .B1(new_n766), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n665), .A2(new_n488), .ZN(new_n775));
  INV_X1    g589(.A(new_n726), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n776), .A2(new_n683), .A3(new_n310), .A4(new_n419), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n778), .A2(new_n412), .A3(new_n751), .ZN(new_n779));
  OR2_X1    g593(.A1(new_n779), .A2(KEYINPUT120), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(KEYINPUT120), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n774), .A2(new_n726), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  AND2_X1   g596(.A1(new_n758), .A2(new_n777), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(new_n720), .ZN(new_n784));
  INV_X1    g598(.A(new_n771), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n667), .A2(new_n312), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n785), .A2(KEYINPUT50), .A3(new_n684), .A4(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n758), .A2(new_n418), .A3(new_n770), .A4(new_n684), .ZN(new_n789));
  INV_X1    g603(.A(new_n786), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n788), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n782), .A2(KEYINPUT51), .A3(new_n784), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n780), .A2(new_n781), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n795), .A2(new_n796), .A3(new_n773), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n726), .A3(new_n785), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n794), .A2(new_n784), .A3(new_n792), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT51), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n684), .A2(new_n364), .ZN(new_n802));
  OAI211_X1 g616(.A(G952), .B(new_n349), .C1(new_n771), .C2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n778), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n803), .B1(new_n610), .B2(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n793), .A2(new_n801), .A3(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n653), .A2(new_n657), .ZN(new_n807));
  AOI211_X1 g621(.A(new_n676), .B(new_n802), .C1(new_n716), .C2(new_n719), .ZN(new_n808));
  OAI21_X1  g622(.A(KEYINPUT118), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n600), .A2(new_n650), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n665), .A3(new_n654), .A4(new_n693), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(KEYINPUT52), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT118), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n721), .A2(new_n658), .A3(new_n813), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n809), .A2(new_n678), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n721), .A2(new_n658), .A3(new_n678), .A4(new_n811), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT52), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n643), .A2(new_n597), .A3(new_n710), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n452), .A2(new_n448), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(KEYINPUT116), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n412), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n612), .B1(new_n611), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n601), .A2(new_n617), .A3(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n685), .A2(new_n825), .A3(new_n688), .A4(new_n691), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n820), .A2(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n600), .A2(new_n650), .A3(new_n776), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n611), .B1(new_n716), .B2(new_n719), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n655), .A2(new_n628), .A3(new_n822), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n728), .A2(new_n730), .A3(new_n733), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n827), .A2(KEYINPUT53), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n819), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(KEYINPUT119), .B(KEYINPUT54), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n721), .A2(new_n658), .A3(new_n678), .ZN(new_n839));
  AOI22_X1  g653(.A1(new_n839), .A2(new_n812), .B1(new_n816), .B2(new_n817), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n643), .A2(new_n597), .A3(new_n710), .ZN(new_n841));
  AND4_X1   g655(.A1(new_n685), .A2(new_n825), .A3(new_n688), .A4(new_n691), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n841), .A2(new_n842), .A3(new_n831), .A4(new_n832), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n838), .B1(new_n840), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n835), .A2(new_n837), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n840), .A2(new_n838), .A3(new_n843), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n843), .A2(KEYINPUT117), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n843), .A2(KEYINPUT117), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n819), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n847), .B1(new_n850), .B2(new_n838), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n806), .B(new_n845), .C1(new_n846), .C2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(new_n725), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n783), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g668(.A(new_n854), .B(KEYINPUT48), .Z(new_n855));
  OAI22_X1  g669(.A1(new_n852), .A2(new_n855), .B1(G952), .B2(G953), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n667), .A2(new_n412), .A3(new_n609), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT49), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n857), .B1(new_n858), .B2(new_n772), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n858), .B2(new_n772), .ZN(new_n860));
  INV_X1    g674(.A(new_n310), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n312), .A3(new_n861), .A4(new_n775), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n856), .A2(new_n862), .ZN(G75));
  AOI21_X1  g677(.A(new_n293), .B1(new_n835), .B2(new_n844), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT56), .B1(new_n864), .B2(G210), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n343), .A2(new_n345), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(new_n351), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT55), .Z(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n865), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n865), .A2(new_n869), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n349), .A2(G952), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT121), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n870), .A2(new_n871), .A3(new_n873), .ZN(G51));
  NAND2_X1  g688(.A1(new_n845), .A2(KEYINPUT122), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n835), .A2(new_n844), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n836), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n835), .A2(new_n844), .A3(new_n878), .A4(new_n837), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n875), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n739), .B(KEYINPUT57), .Z(new_n881));
  NAND2_X1  g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n301), .ZN(new_n883));
  INV_X1    g697(.A(new_n738), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n864), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n872), .B1(new_n883), .B2(new_n885), .ZN(G54));
  NAND2_X1  g700(.A1(new_n394), .A2(new_n401), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n844), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n833), .B1(new_n815), .B2(new_n818), .ZN(new_n890));
  OAI211_X1 g704(.A(KEYINPUT58), .B(G902), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(G475), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n888), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT123), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n872), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n864), .A2(KEYINPUT58), .A3(G475), .A4(new_n887), .ZN(new_n896));
  OAI211_X1 g710(.A(KEYINPUT123), .B(new_n888), .C1(new_n891), .C2(new_n892), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G60));
  NAND2_X1  g712(.A1(new_n606), .A2(new_n607), .ZN(new_n899));
  NAND2_X1  g713(.A1(G478), .A2(G902), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(KEYINPUT59), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n880), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n845), .B1(new_n851), .B2(new_n846), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n899), .B1(new_n904), .B2(new_n901), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n903), .A2(new_n905), .A3(new_n873), .ZN(G63));
  INV_X1    g720(.A(new_n873), .ZN(new_n907));
  NAND2_X1  g721(.A1(G217), .A2(G902), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT60), .Z(new_n909));
  NAND3_X1  g723(.A1(new_n876), .A2(new_n640), .A3(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n876), .A2(new_n909), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n907), .B(new_n910), .C1(new_n911), .C2(new_n478), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(G66));
  INV_X1    g728(.A(G224), .ZN(new_n915));
  OAI21_X1  g729(.A(G953), .B1(new_n414), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n827), .B2(G953), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n866), .B1(G898), .B2(new_n349), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n917), .B(new_n918), .ZN(G69));
  XNOR2_X1  g733(.A(new_n510), .B(new_n397), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n277), .A2(G900), .A3(G953), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n768), .B1(new_n760), .B2(new_n762), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n809), .A2(new_n814), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n678), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n747), .A2(new_n693), .A3(new_n853), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n832), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n923), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  OAI211_X1 g742(.A(new_n921), .B(new_n922), .C1(new_n928), .C2(G953), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n924), .A2(new_n673), .A3(new_n678), .ZN(new_n930));
  XNOR2_X1  g744(.A(KEYINPUT124), .B(KEYINPUT62), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n923), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  AND2_X1   g746(.A1(new_n591), .A2(new_n311), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n611), .A2(new_n823), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n933), .A2(new_n670), .A3(new_n726), .A4(new_n934), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT125), .Z(new_n936));
  AND2_X1   g750(.A1(KEYINPUT124), .A2(KEYINPUT62), .ZN(new_n937));
  OR2_X1    g751(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n932), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n920), .B1(new_n939), .B2(G953), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n277), .A2(new_n649), .A3(new_n349), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n929), .B1(new_n940), .B2(new_n941), .ZN(G72));
  XNOR2_X1  g756(.A(new_n576), .B(KEYINPUT126), .ZN(new_n943));
  INV_X1    g757(.A(new_n827), .ZN(new_n944));
  NOR4_X1   g758(.A1(new_n923), .A2(new_n927), .A3(new_n925), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(G472), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT63), .Z(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n943), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n661), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(new_n576), .A3(new_n947), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT127), .Z(new_n952));
  OAI21_X1  g766(.A(new_n949), .B1(new_n851), .B2(new_n952), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n932), .A2(new_n827), .A3(new_n936), .A4(new_n938), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n950), .B1(new_n954), .B2(new_n947), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n953), .A2(new_n955), .A3(new_n872), .ZN(G57));
endmodule


