

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589;

  XNOR2_X2 U323 ( .A(n458), .B(KEYINPUT122), .ZN(n571) );
  XOR2_X1 U324 ( .A(n374), .B(n349), .Z(n565) );
  XNOR2_X1 U325 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U326 ( .A(n293), .B(n292), .ZN(n398) );
  NOR2_X1 U327 ( .A1(n440), .A2(n514), .ZN(n574) );
  XNOR2_X1 U328 ( .A(n565), .B(n350), .ZN(n549) );
  NOR2_X1 U329 ( .A1(n527), .A2(n526), .ZN(n528) );
  XOR2_X1 U330 ( .A(KEYINPUT112), .B(n533), .Z(n291) );
  INV_X1 U331 ( .A(G106GAT), .ZN(n342) );
  XNOR2_X1 U332 ( .A(n343), .B(n342), .ZN(n345) );
  XNOR2_X1 U333 ( .A(KEYINPUT47), .B(KEYINPUT116), .ZN(n391) );
  XNOR2_X1 U334 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U335 ( .A(n345), .B(n344), .ZN(n361) );
  INV_X1 U336 ( .A(KEYINPUT48), .ZN(n395) );
  XNOR2_X1 U337 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U338 ( .A(n395), .B(KEYINPUT64), .ZN(n396) );
  XNOR2_X1 U339 ( .A(n365), .B(n364), .ZN(n366) );
  AND2_X1 U340 ( .A1(n457), .A2(n519), .ZN(n458) );
  XNOR2_X1 U341 ( .A(n397), .B(n396), .ZN(n556) );
  XNOR2_X1 U342 ( .A(n367), .B(n366), .ZN(n579) );
  XOR2_X1 U343 ( .A(n456), .B(n455), .Z(n519) );
  XNOR2_X1 U344 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U345 ( .A(n462), .B(n461), .ZN(G1349GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT21), .B(G204GAT), .Z(n293) );
  XNOR2_X1 U347 ( .A(G197GAT), .B(G211GAT), .ZN(n292) );
  XOR2_X1 U348 ( .A(KEYINPUT2), .B(KEYINPUT91), .Z(n295) );
  XNOR2_X1 U349 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n294) );
  XNOR2_X1 U350 ( .A(n295), .B(n294), .ZN(n425) );
  XNOR2_X1 U351 ( .A(n398), .B(n425), .ZN(n309) );
  XOR2_X1 U352 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n297) );
  XNOR2_X1 U353 ( .A(G106GAT), .B(KEYINPUT24), .ZN(n296) );
  XNOR2_X1 U354 ( .A(n297), .B(n296), .ZN(n301) );
  XOR2_X1 U355 ( .A(KEYINPUT78), .B(G162GAT), .Z(n346) );
  XOR2_X1 U356 ( .A(G218GAT), .B(n346), .Z(n299) );
  XOR2_X1 U357 ( .A(G22GAT), .B(G141GAT), .Z(n377) );
  XNOR2_X1 U358 ( .A(G50GAT), .B(n377), .ZN(n298) );
  XNOR2_X1 U359 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U360 ( .A(n301), .B(n300), .Z(n303) );
  NAND2_X1 U361 ( .A1(G228GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U362 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U363 ( .A(n304), .B(KEYINPUT92), .Z(n307) );
  XNOR2_X1 U364 ( .A(G78GAT), .B(KEYINPUT74), .ZN(n305) );
  XNOR2_X1 U365 ( .A(n305), .B(G148GAT), .ZN(n358) );
  XNOR2_X1 U366 ( .A(n358), .B(KEYINPUT90), .ZN(n306) );
  XNOR2_X1 U367 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n475) );
  XNOR2_X1 U369 ( .A(KEYINPUT121), .B(KEYINPUT54), .ZN(n415) );
  XOR2_X1 U370 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n311) );
  XNOR2_X1 U371 ( .A(G78GAT), .B(G64GAT), .ZN(n310) );
  XNOR2_X1 U372 ( .A(n311), .B(n310), .ZN(n325) );
  XOR2_X1 U373 ( .A(KEYINPUT13), .B(G57GAT), .Z(n352) );
  XOR2_X1 U374 ( .A(n352), .B(G211GAT), .Z(n314) );
  XNOR2_X1 U375 ( .A(G1GAT), .B(KEYINPUT71), .ZN(n312) );
  XNOR2_X1 U376 ( .A(n312), .B(G15GAT), .ZN(n379) );
  XNOR2_X1 U377 ( .A(n379), .B(G22GAT), .ZN(n313) );
  XNOR2_X1 U378 ( .A(n314), .B(n313), .ZN(n318) );
  XOR2_X1 U379 ( .A(G127GAT), .B(G155GAT), .Z(n316) );
  NAND2_X1 U380 ( .A1(G231GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U381 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U382 ( .A(n318), .B(n317), .Z(n323) );
  XOR2_X1 U383 ( .A(KEYINPUT12), .B(KEYINPUT84), .Z(n320) );
  XNOR2_X1 U384 ( .A(G183GAT), .B(G71GAT), .ZN(n319) );
  XNOR2_X1 U385 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U386 ( .A(G8GAT), .B(n321), .ZN(n322) );
  XNOR2_X1 U387 ( .A(n323), .B(n322), .ZN(n324) );
  XOR2_X1 U388 ( .A(n325), .B(n324), .Z(n495) );
  XOR2_X1 U389 ( .A(G43GAT), .B(G29GAT), .Z(n327) );
  XNOR2_X1 U390 ( .A(KEYINPUT70), .B(G50GAT), .ZN(n326) );
  XNOR2_X1 U391 ( .A(n327), .B(n326), .ZN(n329) );
  INV_X1 U392 ( .A(KEYINPUT7), .ZN(n328) );
  XNOR2_X1 U393 ( .A(n329), .B(n328), .ZN(n331) );
  XNOR2_X1 U394 ( .A(G36GAT), .B(KEYINPUT8), .ZN(n330) );
  XNOR2_X1 U395 ( .A(n331), .B(n330), .ZN(n374) );
  XOR2_X1 U396 ( .A(KEYINPUT79), .B(KEYINPUT81), .Z(n333) );
  XNOR2_X1 U397 ( .A(KEYINPUT11), .B(KEYINPUT65), .ZN(n332) );
  XNOR2_X1 U398 ( .A(n333), .B(n332), .ZN(n335) );
  INV_X1 U399 ( .A(KEYINPUT10), .ZN(n334) );
  XNOR2_X1 U400 ( .A(n335), .B(n334), .ZN(n337) );
  XOR2_X1 U401 ( .A(G190GAT), .B(G218GAT), .Z(n405) );
  XNOR2_X1 U402 ( .A(n405), .B(KEYINPUT80), .ZN(n336) );
  XNOR2_X1 U403 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U404 ( .A(G134GAT), .B(KEYINPUT82), .Z(n430) );
  XOR2_X1 U405 ( .A(n430), .B(KEYINPUT9), .Z(n339) );
  NAND2_X1 U406 ( .A1(G232GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U407 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U408 ( .A(n341), .B(n340), .ZN(n348) );
  XNOR2_X1 U409 ( .A(G99GAT), .B(G92GAT), .ZN(n343) );
  XOR2_X1 U410 ( .A(KEYINPUT75), .B(G85GAT), .Z(n344) );
  XOR2_X1 U411 ( .A(n361), .B(n346), .Z(n347) );
  XNOR2_X1 U412 ( .A(n348), .B(n347), .ZN(n349) );
  INV_X1 U413 ( .A(KEYINPUT83), .ZN(n350) );
  XOR2_X1 U414 ( .A(KEYINPUT36), .B(n549), .Z(n586) );
  NOR2_X1 U415 ( .A1(n495), .A2(n586), .ZN(n351) );
  XNOR2_X1 U416 ( .A(KEYINPUT45), .B(n351), .ZN(n384) );
  XOR2_X1 U417 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n354) );
  XOR2_X1 U418 ( .A(G176GAT), .B(G64GAT), .Z(n401) );
  XNOR2_X1 U419 ( .A(n352), .B(n401), .ZN(n353) );
  XNOR2_X1 U420 ( .A(n354), .B(n353), .ZN(n360) );
  NAND2_X1 U421 ( .A1(G230GAT), .A2(G233GAT), .ZN(n356) );
  INV_X1 U422 ( .A(KEYINPUT33), .ZN(n355) );
  XOR2_X1 U423 ( .A(n360), .B(n359), .Z(n367) );
  XOR2_X1 U424 ( .A(G71GAT), .B(G120GAT), .Z(n444) );
  XNOR2_X1 U425 ( .A(n444), .B(n361), .ZN(n365) );
  XOR2_X1 U426 ( .A(KEYINPUT31), .B(KEYINPUT76), .Z(n363) );
  XNOR2_X1 U427 ( .A(G204GAT), .B(KEYINPUT77), .ZN(n362) );
  XOR2_X1 U428 ( .A(n363), .B(n362), .Z(n364) );
  XOR2_X1 U429 ( .A(KEYINPUT30), .B(KEYINPUT69), .Z(n369) );
  NAND2_X1 U430 ( .A1(G229GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U431 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U432 ( .A(n370), .B(G197GAT), .Z(n376) );
  XOR2_X1 U433 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n372) );
  XNOR2_X1 U434 ( .A(G113GAT), .B(KEYINPUT67), .ZN(n371) );
  XNOR2_X1 U435 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U437 ( .A(n376), .B(n375), .ZN(n378) );
  XNOR2_X1 U438 ( .A(n378), .B(n377), .ZN(n381) );
  XOR2_X1 U439 ( .A(G169GAT), .B(G8GAT), .Z(n411) );
  XOR2_X1 U440 ( .A(n379), .B(n411), .Z(n380) );
  XNOR2_X1 U441 ( .A(n381), .B(n380), .ZN(n575) );
  XNOR2_X1 U442 ( .A(KEYINPUT72), .B(n575), .ZN(n568) );
  INV_X1 U443 ( .A(n568), .ZN(n382) );
  AND2_X1 U444 ( .A1(n579), .A2(n382), .ZN(n383) );
  AND2_X1 U445 ( .A1(n384), .A2(n383), .ZN(n385) );
  XNOR2_X1 U446 ( .A(n385), .B(KEYINPUT117), .ZN(n394) );
  XNOR2_X1 U447 ( .A(n579), .B(KEYINPUT41), .ZN(n560) );
  AND2_X1 U448 ( .A1(n575), .A2(n560), .ZN(n387) );
  INV_X1 U449 ( .A(KEYINPUT46), .ZN(n386) );
  XNOR2_X1 U450 ( .A(n387), .B(n386), .ZN(n388) );
  AND2_X1 U451 ( .A1(n388), .A2(n495), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n389), .B(KEYINPUT115), .ZN(n390) );
  NOR2_X1 U453 ( .A1(n565), .A2(n390), .ZN(n392) );
  NAND2_X1 U454 ( .A1(n394), .A2(n393), .ZN(n397) );
  XOR2_X1 U455 ( .A(KEYINPUT96), .B(n398), .Z(n400) );
  NAND2_X1 U456 ( .A1(G226GAT), .A2(G233GAT), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n402) );
  XOR2_X1 U458 ( .A(n402), .B(n401), .Z(n404) );
  XNOR2_X1 U459 ( .A(G36GAT), .B(G92GAT), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n406) );
  XOR2_X1 U461 ( .A(n406), .B(n405), .Z(n413) );
  XNOR2_X1 U462 ( .A(KEYINPUT89), .B(KEYINPUT17), .ZN(n407) );
  XNOR2_X1 U463 ( .A(n407), .B(KEYINPUT88), .ZN(n408) );
  XOR2_X1 U464 ( .A(n408), .B(KEYINPUT19), .Z(n410) );
  XNOR2_X1 U465 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n410), .B(n409), .ZN(n452) );
  XNOR2_X1 U467 ( .A(n411), .B(n452), .ZN(n412) );
  XNOR2_X1 U468 ( .A(n413), .B(n412), .ZN(n532) );
  NOR2_X1 U469 ( .A1(n556), .A2(n532), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n415), .B(n414), .ZN(n440) );
  XOR2_X1 U471 ( .A(G127GAT), .B(KEYINPUT0), .Z(n417) );
  XNOR2_X1 U472 ( .A(G113GAT), .B(KEYINPUT86), .ZN(n416) );
  XNOR2_X1 U473 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U474 ( .A(KEYINPUT85), .B(n418), .ZN(n455) );
  INV_X1 U475 ( .A(n455), .ZN(n439) );
  XOR2_X1 U476 ( .A(KEYINPUT93), .B(KEYINPUT95), .Z(n420) );
  XNOR2_X1 U477 ( .A(G120GAT), .B(G148GAT), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U479 ( .A(KEYINPUT94), .B(KEYINPUT4), .Z(n422) );
  XNOR2_X1 U480 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n421) );
  XNOR2_X1 U481 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U482 ( .A(n424), .B(n423), .Z(n437) );
  XOR2_X1 U483 ( .A(n425), .B(KEYINPUT5), .Z(n427) );
  NAND2_X1 U484 ( .A1(G225GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n435) );
  XOR2_X1 U486 ( .A(G57GAT), .B(G162GAT), .Z(n429) );
  XNOR2_X1 U487 ( .A(G1GAT), .B(G141GAT), .ZN(n428) );
  XNOR2_X1 U488 ( .A(n429), .B(n428), .ZN(n431) );
  XOR2_X1 U489 ( .A(n431), .B(n430), .Z(n433) );
  XNOR2_X1 U490 ( .A(G29GAT), .B(G85GAT), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U494 ( .A(n439), .B(n438), .Z(n529) );
  INV_X1 U495 ( .A(n529), .ZN(n514) );
  NAND2_X1 U496 ( .A1(n475), .A2(n574), .ZN(n441) );
  XNOR2_X1 U497 ( .A(KEYINPUT55), .B(n441), .ZN(n457) );
  XOR2_X1 U498 ( .A(G190GAT), .B(G134GAT), .Z(n443) );
  XNOR2_X1 U499 ( .A(G43GAT), .B(G99GAT), .ZN(n442) );
  XNOR2_X1 U500 ( .A(n443), .B(n442), .ZN(n445) );
  XOR2_X1 U501 ( .A(n445), .B(n444), .Z(n447) );
  XNOR2_X1 U502 ( .A(G169GAT), .B(G15GAT), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U504 ( .A(KEYINPUT20), .B(KEYINPUT87), .Z(n449) );
  NAND2_X1 U505 ( .A1(G227GAT), .A2(G233GAT), .ZN(n448) );
  XNOR2_X1 U506 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U507 ( .A(n451), .B(n450), .Z(n454) );
  XNOR2_X1 U508 ( .A(n452), .B(G176GAT), .ZN(n453) );
  XNOR2_X1 U509 ( .A(n454), .B(n453), .ZN(n456) );
  NAND2_X1 U510 ( .A1(n571), .A2(n560), .ZN(n462) );
  XOR2_X1 U511 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n460) );
  XNOR2_X1 U512 ( .A(G176GAT), .B(KEYINPUT124), .ZN(n459) );
  NAND2_X1 U513 ( .A1(n571), .A2(n549), .ZN(n466) );
  XNOR2_X1 U514 ( .A(G190GAT), .B(KEYINPUT126), .ZN(n463) );
  XNOR2_X1 U515 ( .A(n463), .B(KEYINPUT125), .ZN(n464) );
  XOR2_X1 U516 ( .A(KEYINPUT58), .B(n464), .Z(n465) );
  XNOR2_X1 U517 ( .A(n466), .B(n465), .ZN(G1351GAT) );
  XOR2_X1 U518 ( .A(KEYINPUT34), .B(KEYINPUT103), .Z(n487) );
  NOR2_X1 U519 ( .A1(n495), .A2(n549), .ZN(n467) );
  XNOR2_X1 U520 ( .A(KEYINPUT16), .B(n467), .ZN(n484) );
  XNOR2_X1 U521 ( .A(n475), .B(KEYINPUT28), .ZN(n468) );
  XNOR2_X1 U522 ( .A(n468), .B(KEYINPUT66), .ZN(n538) );
  XNOR2_X1 U523 ( .A(n532), .B(KEYINPUT97), .ZN(n469) );
  XNOR2_X1 U524 ( .A(n469), .B(KEYINPUT27), .ZN(n478) );
  NAND2_X1 U525 ( .A1(n478), .A2(n514), .ZN(n470) );
  XOR2_X1 U526 ( .A(KEYINPUT98), .B(n470), .Z(n554) );
  NAND2_X1 U527 ( .A1(n538), .A2(n554), .ZN(n542) );
  XNOR2_X1 U528 ( .A(n542), .B(KEYINPUT99), .ZN(n471) );
  INV_X1 U529 ( .A(n519), .ZN(n541) );
  NAND2_X1 U530 ( .A1(n471), .A2(n541), .ZN(n483) );
  INV_X1 U531 ( .A(n532), .ZN(n517) );
  NAND2_X1 U532 ( .A1(n519), .A2(n517), .ZN(n472) );
  NAND2_X1 U533 ( .A1(n472), .A2(n475), .ZN(n473) );
  XNOR2_X1 U534 ( .A(n473), .B(KEYINPUT25), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n474), .B(KEYINPUT101), .ZN(n480) );
  NOR2_X1 U536 ( .A1(n475), .A2(n519), .ZN(n477) );
  XNOR2_X1 U537 ( .A(KEYINPUT26), .B(KEYINPUT100), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(n573) );
  NAND2_X1 U539 ( .A1(n478), .A2(n573), .ZN(n479) );
  NAND2_X1 U540 ( .A1(n480), .A2(n479), .ZN(n481) );
  NAND2_X1 U541 ( .A1(n529), .A2(n481), .ZN(n482) );
  NAND2_X1 U542 ( .A1(n483), .A2(n482), .ZN(n496) );
  NAND2_X1 U543 ( .A1(n484), .A2(n496), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n485), .B(KEYINPUT102), .ZN(n513) );
  NAND2_X1 U545 ( .A1(n579), .A2(n568), .ZN(n500) );
  NOR2_X1 U546 ( .A1(n513), .A2(n500), .ZN(n493) );
  NAND2_X1 U547 ( .A1(n493), .A2(n514), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n488), .ZN(G1324GAT) );
  NAND2_X1 U550 ( .A1(n517), .A2(n493), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n489), .B(KEYINPUT104), .ZN(n490) );
  XNOR2_X1 U552 ( .A(G8GAT), .B(n490), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT35), .Z(n492) );
  NAND2_X1 U554 ( .A1(n493), .A2(n519), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(G1326GAT) );
  INV_X1 U556 ( .A(n538), .ZN(n521) );
  NAND2_X1 U557 ( .A1(n521), .A2(n493), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n494), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT106), .Z(n503) );
  XNOR2_X1 U560 ( .A(KEYINPUT37), .B(KEYINPUT105), .ZN(n499) );
  INV_X1 U561 ( .A(n495), .ZN(n583) );
  NOR2_X1 U562 ( .A1(n586), .A2(n583), .ZN(n497) );
  NAND2_X1 U563 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n499), .B(n498), .ZN(n527) );
  NOR2_X1 U565 ( .A1(n500), .A2(n527), .ZN(n501) );
  XNOR2_X1 U566 ( .A(n501), .B(KEYINPUT38), .ZN(n509) );
  NAND2_X1 U567 ( .A1(n509), .A2(n514), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(n505) );
  XOR2_X1 U569 ( .A(KEYINPUT39), .B(KEYINPUT107), .Z(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(G1328GAT) );
  NAND2_X1 U571 ( .A1(n509), .A2(n517), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n506), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U573 ( .A1(n509), .A2(n519), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n507), .B(KEYINPUT40), .ZN(n508) );
  XNOR2_X1 U575 ( .A(G43GAT), .B(n508), .ZN(G1330GAT) );
  NAND2_X1 U576 ( .A1(n509), .A2(n521), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n510), .B(KEYINPUT108), .ZN(n511) );
  XNOR2_X1 U578 ( .A(G50GAT), .B(n511), .ZN(G1331GAT) );
  XNOR2_X1 U579 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n516) );
  INV_X1 U580 ( .A(n575), .ZN(n512) );
  NAND2_X1 U581 ( .A1(n512), .A2(n560), .ZN(n526) );
  NOR2_X1 U582 ( .A1(n513), .A2(n526), .ZN(n522) );
  NAND2_X1 U583 ( .A1(n522), .A2(n514), .ZN(n515) );
  XNOR2_X1 U584 ( .A(n516), .B(n515), .ZN(G1332GAT) );
  NAND2_X1 U585 ( .A1(n517), .A2(n522), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n518), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U587 ( .A1(n519), .A2(n522), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n520), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U589 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n524) );
  NAND2_X1 U590 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U592 ( .A(G78GAT), .B(n525), .Z(G1335GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT110), .B(n528), .Z(n537) );
  NOR2_X1 U594 ( .A1(n529), .A2(n537), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n530), .B(KEYINPUT111), .ZN(n531) );
  XNOR2_X1 U596 ( .A(G85GAT), .B(n531), .ZN(G1336GAT) );
  NOR2_X1 U597 ( .A1(n532), .A2(n537), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G92GAT), .B(n291), .ZN(G1337GAT) );
  NOR2_X1 U599 ( .A1(n541), .A2(n537), .ZN(n534) );
  XOR2_X1 U600 ( .A(G99GAT), .B(n534), .Z(G1338GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n536) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(KEYINPUT114), .ZN(n535) );
  XNOR2_X1 U603 ( .A(n536), .B(n535), .ZN(n540) );
  NOR2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U605 ( .A(n540), .B(n539), .Z(G1339GAT) );
  OR2_X1 U606 ( .A1(n542), .A2(n541), .ZN(n543) );
  NOR2_X1 U607 ( .A1(n556), .A2(n543), .ZN(n550) );
  NAND2_X1 U608 ( .A1(n550), .A2(n568), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G113GAT), .B(n544), .ZN(G1340GAT) );
  XOR2_X1 U610 ( .A(G120GAT), .B(KEYINPUT49), .Z(n546) );
  NAND2_X1 U611 ( .A1(n550), .A2(n560), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1341GAT) );
  NAND2_X1 U613 ( .A1(n583), .A2(n550), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n547), .B(KEYINPUT50), .ZN(n548) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT51), .B(KEYINPUT118), .Z(n552) );
  NAND2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(G134GAT), .B(n553), .ZN(G1343GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n558) );
  NAND2_X1 U621 ( .A1(n573), .A2(n554), .ZN(n555) );
  NOR2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n566), .A2(n575), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G141GAT), .B(n559), .ZN(G1344GAT) );
  XOR2_X1 U626 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n562) );
  NAND2_X1 U627 ( .A1(n566), .A2(n560), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G148GAT), .B(n563), .ZN(G1345GAT) );
  NAND2_X1 U630 ( .A1(n583), .A2(n566), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U632 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n567), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U634 ( .A(G169GAT), .B(KEYINPUT123), .Z(n570) );
  NAND2_X1 U635 ( .A1(n571), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(G1348GAT) );
  NAND2_X1 U637 ( .A1(n571), .A2(n583), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n577) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n585) );
  INV_X1 U641 ( .A(n585), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n582), .A2(n575), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  XOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .Z(n581) );
  OR2_X1 U646 ( .A1(n585), .A2(n579), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n584), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U651 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U653 ( .A(G218GAT), .B(n589), .ZN(G1355GAT) );
endmodule

