

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U553 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X2 U554 ( .A1(n543), .A2(G543), .ZN(n541) );
  INV_X2 U555 ( .A(n724), .ZN(n709) );
  XNOR2_X2 U556 ( .A(n528), .B(KEYINPUT64), .ZN(n666) );
  AND2_X1 U557 ( .A1(n526), .A2(n525), .ZN(n674) );
  AND2_X2 U558 ( .A1(G2105), .A2(G2104), .ZN(n888) );
  NAND2_X1 U559 ( .A1(n888), .A2(G113), .ZN(n519) );
  XOR2_X1 U560 ( .A(KEYINPUT65), .B(n519), .Z(n522) );
  NOR2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XOR2_X1 U562 ( .A(KEYINPUT17), .B(n520), .Z(n530) );
  NAND2_X1 U563 ( .A1(n530), .A2(G137), .ZN(n521) );
  NAND2_X1 U564 ( .A1(n522), .A2(n521), .ZN(n524) );
  INV_X1 U565 ( .A(KEYINPUT66), .ZN(n523) );
  XNOR2_X1 U566 ( .A(n524), .B(n523), .ZN(n526) );
  INV_X1 U567 ( .A(G2105), .ZN(n527) );
  NOR2_X1 U568 ( .A1(G2104), .A2(n527), .ZN(n887) );
  NAND2_X1 U569 ( .A1(n887), .A2(G125), .ZN(n525) );
  AND2_X1 U570 ( .A1(G2104), .A2(n527), .ZN(n528) );
  NAND2_X1 U571 ( .A1(G101), .A2(n666), .ZN(n529) );
  XOR2_X1 U572 ( .A(KEYINPUT23), .B(n529), .Z(n673) );
  AND2_X1 U573 ( .A1(n674), .A2(n673), .ZN(G160) );
  AND2_X1 U574 ( .A1(G452), .A2(G94), .ZN(G173) );
  BUF_X1 U575 ( .A(n530), .Z(n893) );
  NAND2_X1 U576 ( .A1(G135), .A2(n893), .ZN(n531) );
  XNOR2_X1 U577 ( .A(n531), .B(KEYINPUT78), .ZN(n538) );
  NAND2_X1 U578 ( .A1(n888), .A2(G111), .ZN(n533) );
  NAND2_X1 U579 ( .A1(G99), .A2(n666), .ZN(n532) );
  NAND2_X1 U580 ( .A1(n533), .A2(n532), .ZN(n536) );
  NAND2_X1 U581 ( .A1(n887), .A2(G123), .ZN(n534) );
  XOR2_X1 U582 ( .A(KEYINPUT18), .B(n534), .Z(n535) );
  NOR2_X1 U583 ( .A1(n536), .A2(n535), .ZN(n537) );
  NAND2_X1 U584 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U585 ( .A(KEYINPUT79), .B(n539), .Z(n994) );
  XNOR2_X1 U586 ( .A(G2096), .B(n994), .ZN(n540) );
  OR2_X1 U587 ( .A1(G2100), .A2(n540), .ZN(G156) );
  INV_X1 U588 ( .A(G108), .ZN(G238) );
  INV_X1 U589 ( .A(G120), .ZN(G236) );
  INV_X1 U590 ( .A(G69), .ZN(G235) );
  INV_X1 U591 ( .A(G132), .ZN(G219) );
  INV_X1 U592 ( .A(G82), .ZN(G220) );
  XNOR2_X1 U593 ( .A(KEYINPUT67), .B(G651), .ZN(n543) );
  XOR2_X2 U594 ( .A(KEYINPUT1), .B(n541), .Z(n634) );
  NAND2_X1 U595 ( .A1(G64), .A2(n634), .ZN(n542) );
  XNOR2_X1 U596 ( .A(KEYINPUT69), .B(n542), .ZN(n551) );
  NOR2_X1 U597 ( .A1(G651), .A2(G543), .ZN(n633) );
  NAND2_X1 U598 ( .A1(G90), .A2(n633), .ZN(n545) );
  XOR2_X1 U599 ( .A(G543), .B(KEYINPUT0), .Z(n611) );
  NOR2_X4 U600 ( .A1(n611), .A2(n543), .ZN(n638) );
  NAND2_X1 U601 ( .A1(G77), .A2(n638), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U603 ( .A(n546), .B(KEYINPUT70), .ZN(n547) );
  XNOR2_X1 U604 ( .A(n547), .B(KEYINPUT9), .ZN(n549) );
  NOR2_X2 U605 ( .A1(G651), .A2(n611), .ZN(n637) );
  NAND2_X1 U606 ( .A1(n637), .A2(G52), .ZN(n548) );
  NAND2_X1 U607 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U608 ( .A1(n551), .A2(n550), .ZN(G171) );
  NAND2_X1 U609 ( .A1(n637), .A2(G51), .ZN(n553) );
  NAND2_X1 U610 ( .A1(G63), .A2(n634), .ZN(n552) );
  NAND2_X1 U611 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U612 ( .A(KEYINPUT6), .B(n554), .ZN(n560) );
  NAND2_X1 U613 ( .A1(n633), .A2(G89), .ZN(n555) );
  XNOR2_X1 U614 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G76), .A2(n638), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U617 ( .A(n558), .B(KEYINPUT5), .Z(n559) );
  NOR2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U619 ( .A(KEYINPUT75), .B(n561), .Z(n562) );
  XOR2_X1 U620 ( .A(KEYINPUT7), .B(n562), .Z(G168) );
  XOR2_X1 U621 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U622 ( .A1(G7), .A2(G661), .ZN(n563) );
  XNOR2_X1 U623 ( .A(n563), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U624 ( .A(G223), .ZN(n832) );
  NAND2_X1 U625 ( .A1(n832), .A2(G567), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  NAND2_X1 U627 ( .A1(n634), .A2(G56), .ZN(n565) );
  XOR2_X1 U628 ( .A(KEYINPUT14), .B(n565), .Z(n571) );
  NAND2_X1 U629 ( .A1(n633), .A2(G81), .ZN(n566) );
  XNOR2_X1 U630 ( .A(n566), .B(KEYINPUT12), .ZN(n568) );
  NAND2_X1 U631 ( .A1(G68), .A2(n638), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT13), .B(n569), .Z(n570) );
  NOR2_X1 U634 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n637), .A2(G43), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n573), .A2(n572), .ZN(n941) );
  INV_X1 U637 ( .A(G860), .ZN(n837) );
  OR2_X1 U638 ( .A1(n941), .A2(n837), .ZN(G153) );
  INV_X1 U639 ( .A(G171), .ZN(G301) );
  NAND2_X1 U640 ( .A1(G92), .A2(n633), .ZN(n575) );
  NAND2_X1 U641 ( .A1(G54), .A2(n637), .ZN(n574) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U643 ( .A1(G79), .A2(n638), .ZN(n576) );
  XNOR2_X1 U644 ( .A(n576), .B(KEYINPUT73), .ZN(n577) );
  NOR2_X1 U645 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U646 ( .A1(G66), .A2(n634), .ZN(n579) );
  NAND2_X1 U647 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U648 ( .A(KEYINPUT15), .B(n581), .Z(n582) );
  XNOR2_X1 U649 ( .A(KEYINPUT74), .B(n582), .ZN(n686) );
  BUF_X1 U650 ( .A(n686), .Z(n918) );
  NOR2_X1 U651 ( .A1(n918), .A2(G868), .ZN(n584) );
  INV_X1 U652 ( .A(G868), .ZN(n649) );
  NOR2_X1 U653 ( .A1(n649), .A2(G301), .ZN(n583) );
  NOR2_X1 U654 ( .A1(n584), .A2(n583), .ZN(G284) );
  NAND2_X1 U655 ( .A1(n637), .A2(G53), .ZN(n586) );
  NAND2_X1 U656 ( .A1(G78), .A2(n638), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n590) );
  NAND2_X1 U658 ( .A1(n633), .A2(G91), .ZN(n588) );
  NAND2_X1 U659 ( .A1(G65), .A2(n634), .ZN(n587) );
  NAND2_X1 U660 ( .A1(n588), .A2(n587), .ZN(n589) );
  NOR2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U662 ( .A(n591), .B(KEYINPUT71), .ZN(n919) );
  XNOR2_X1 U663 ( .A(KEYINPUT72), .B(n919), .ZN(G299) );
  NOR2_X1 U664 ( .A1(G286), .A2(n649), .ZN(n592) );
  XNOR2_X1 U665 ( .A(n592), .B(KEYINPUT76), .ZN(n594) );
  NOR2_X1 U666 ( .A1(G299), .A2(G868), .ZN(n593) );
  NOR2_X1 U667 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U668 ( .A1(n837), .A2(G559), .ZN(n595) );
  INV_X1 U669 ( .A(n918), .ZN(n630) );
  NAND2_X1 U670 ( .A1(n595), .A2(n630), .ZN(n596) );
  XNOR2_X1 U671 ( .A(n596), .B(KEYINPUT77), .ZN(n597) );
  XOR2_X1 U672 ( .A(KEYINPUT16), .B(n597), .Z(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n941), .ZN(n600) );
  NAND2_X1 U674 ( .A1(n630), .A2(G868), .ZN(n598) );
  NOR2_X1 U675 ( .A1(G559), .A2(n598), .ZN(n599) );
  NOR2_X1 U676 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U677 ( .A1(G86), .A2(n633), .ZN(n602) );
  NAND2_X1 U678 ( .A1(G48), .A2(n637), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n605) );
  NAND2_X1 U680 ( .A1(n638), .A2(G73), .ZN(n603) );
  XOR2_X1 U681 ( .A(KEYINPUT2), .B(n603), .Z(n604) );
  NOR2_X1 U682 ( .A1(n605), .A2(n604), .ZN(n607) );
  NAND2_X1 U683 ( .A1(G61), .A2(n634), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n607), .A2(n606), .ZN(G305) );
  NAND2_X1 U685 ( .A1(G49), .A2(n637), .ZN(n609) );
  NAND2_X1 U686 ( .A1(G74), .A2(G651), .ZN(n608) );
  NAND2_X1 U687 ( .A1(n609), .A2(n608), .ZN(n610) );
  NOR2_X1 U688 ( .A1(n634), .A2(n610), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G87), .A2(n611), .ZN(n612) );
  XOR2_X1 U690 ( .A(KEYINPUT81), .B(n612), .Z(n613) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(G288) );
  NAND2_X1 U692 ( .A1(n637), .A2(G50), .ZN(n621) );
  NAND2_X1 U693 ( .A1(G62), .A2(n634), .ZN(n616) );
  NAND2_X1 U694 ( .A1(G75), .A2(n638), .ZN(n615) );
  NAND2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U696 ( .A1(n633), .A2(G88), .ZN(n617) );
  XOR2_X1 U697 ( .A(KEYINPUT82), .B(n617), .Z(n618) );
  NOR2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U699 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U700 ( .A(n622), .B(KEYINPUT83), .ZN(G166) );
  NAND2_X1 U701 ( .A1(G85), .A2(n633), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G72), .A2(n638), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U704 ( .A(KEYINPUT68), .B(n625), .Z(n629) );
  NAND2_X1 U705 ( .A1(n634), .A2(G60), .ZN(n627) );
  NAND2_X1 U706 ( .A1(n637), .A2(G47), .ZN(n626) );
  AND2_X1 U707 ( .A1(n627), .A2(n626), .ZN(n628) );
  NAND2_X1 U708 ( .A1(n629), .A2(n628), .ZN(G290) );
  NAND2_X1 U709 ( .A1(n630), .A2(G559), .ZN(n631) );
  XOR2_X1 U710 ( .A(n941), .B(n631), .Z(n836) );
  XNOR2_X1 U711 ( .A(KEYINPUT19), .B(G305), .ZN(n632) );
  XNOR2_X1 U712 ( .A(n632), .B(G288), .ZN(n644) );
  NAND2_X1 U713 ( .A1(n633), .A2(G93), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G67), .A2(n634), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n642) );
  NAND2_X1 U716 ( .A1(n637), .A2(G55), .ZN(n640) );
  NAND2_X1 U717 ( .A1(G80), .A2(n638), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U719 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U720 ( .A(KEYINPUT80), .B(n643), .Z(n838) );
  XOR2_X1 U721 ( .A(n644), .B(n838), .Z(n646) );
  XNOR2_X1 U722 ( .A(G166), .B(G299), .ZN(n645) );
  XNOR2_X1 U723 ( .A(n646), .B(n645), .ZN(n647) );
  XNOR2_X1 U724 ( .A(n647), .B(G290), .ZN(n904) );
  XNOR2_X1 U725 ( .A(n836), .B(n904), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n648), .A2(G868), .ZN(n651) );
  NAND2_X1 U727 ( .A1(n838), .A2(n649), .ZN(n650) );
  NAND2_X1 U728 ( .A1(n651), .A2(n650), .ZN(G295) );
  NAND2_X1 U729 ( .A1(G2078), .A2(G2084), .ZN(n652) );
  XOR2_X1 U730 ( .A(KEYINPUT20), .B(n652), .Z(n653) );
  NAND2_X1 U731 ( .A1(G2090), .A2(n653), .ZN(n654) );
  XNOR2_X1 U732 ( .A(KEYINPUT21), .B(n654), .ZN(n655) );
  NAND2_X1 U733 ( .A1(n655), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U734 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U735 ( .A1(G220), .A2(G219), .ZN(n656) );
  XOR2_X1 U736 ( .A(KEYINPUT22), .B(n656), .Z(n657) );
  NOR2_X1 U737 ( .A1(G218), .A2(n657), .ZN(n658) );
  NAND2_X1 U738 ( .A1(G96), .A2(n658), .ZN(n840) );
  NAND2_X1 U739 ( .A1(n840), .A2(G2106), .ZN(n664) );
  NOR2_X1 U740 ( .A1(G235), .A2(G236), .ZN(n659) );
  XNOR2_X1 U741 ( .A(KEYINPUT84), .B(n659), .ZN(n660) );
  NAND2_X1 U742 ( .A1(n660), .A2(G57), .ZN(n661) );
  NOR2_X1 U743 ( .A1(n661), .A2(G238), .ZN(n662) );
  XNOR2_X1 U744 ( .A(n662), .B(KEYINPUT85), .ZN(n841) );
  NAND2_X1 U745 ( .A1(n841), .A2(G567), .ZN(n663) );
  NAND2_X1 U746 ( .A1(n664), .A2(n663), .ZN(n862) );
  NAND2_X1 U747 ( .A1(G661), .A2(G483), .ZN(n665) );
  NOR2_X1 U748 ( .A1(n862), .A2(n665), .ZN(n835) );
  NAND2_X1 U749 ( .A1(n835), .A2(G36), .ZN(G176) );
  NAND2_X1 U750 ( .A1(n893), .A2(G138), .ZN(n668) );
  NAND2_X1 U751 ( .A1(G102), .A2(n666), .ZN(n667) );
  NAND2_X1 U752 ( .A1(n668), .A2(n667), .ZN(n672) );
  NAND2_X1 U753 ( .A1(G126), .A2(n887), .ZN(n670) );
  NAND2_X1 U754 ( .A1(G114), .A2(n888), .ZN(n669) );
  NAND2_X1 U755 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U756 ( .A1(n672), .A2(n671), .ZN(G164) );
  INV_X1 U757 ( .A(G166), .ZN(G303) );
  NAND2_X1 U758 ( .A1(G1976), .A2(G288), .ZN(n925) );
  AND2_X1 U759 ( .A1(G40), .A2(n673), .ZN(n675) );
  NAND2_X1 U760 ( .A1(n675), .A2(n674), .ZN(n749) );
  XNOR2_X1 U761 ( .A(KEYINPUT91), .B(n749), .ZN(n676) );
  NOR2_X1 U762 ( .A1(G164), .A2(G1384), .ZN(n750) );
  NAND2_X2 U763 ( .A1(n676), .A2(n750), .ZN(n724) );
  NAND2_X1 U764 ( .A1(G8), .A2(n724), .ZN(n797) );
  NAND2_X1 U765 ( .A1(n709), .A2(G2072), .ZN(n677) );
  XOR2_X1 U766 ( .A(KEYINPUT27), .B(n677), .Z(n679) );
  NAND2_X1 U767 ( .A1(G1956), .A2(n724), .ZN(n678) );
  NAND2_X1 U768 ( .A1(n679), .A2(n678), .ZN(n703) );
  NOR2_X1 U769 ( .A1(n919), .A2(n703), .ZN(n680) );
  XNOR2_X1 U770 ( .A(KEYINPUT96), .B(n680), .ZN(n702) );
  AND2_X1 U771 ( .A1(n686), .A2(G1348), .ZN(n683) );
  XNOR2_X1 U772 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n690) );
  INV_X1 U773 ( .A(G1341), .ZN(n681) );
  NAND2_X1 U774 ( .A1(n690), .A2(n681), .ZN(n682) );
  NOR2_X1 U775 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U776 ( .A1(n684), .A2(n709), .ZN(n685) );
  NOR2_X1 U777 ( .A1(n941), .A2(n685), .ZN(n694) );
  NAND2_X1 U778 ( .A1(n686), .A2(G2067), .ZN(n688) );
  NAND2_X1 U779 ( .A1(G1996), .A2(n690), .ZN(n687) );
  NAND2_X1 U780 ( .A1(n688), .A2(n687), .ZN(n689) );
  AND2_X1 U781 ( .A1(n689), .A2(n709), .ZN(n692) );
  NOR2_X1 U782 ( .A1(G1996), .A2(n690), .ZN(n691) );
  NOR2_X1 U783 ( .A1(n692), .A2(n691), .ZN(n693) );
  AND2_X1 U784 ( .A1(n694), .A2(n693), .ZN(n699) );
  NAND2_X1 U785 ( .A1(G1348), .A2(n724), .ZN(n696) );
  NAND2_X1 U786 ( .A1(n709), .A2(G2067), .ZN(n695) );
  NAND2_X1 U787 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U788 ( .A1(n918), .A2(n697), .ZN(n698) );
  XNOR2_X1 U789 ( .A(n700), .B(KEYINPUT95), .ZN(n701) );
  NOR2_X1 U790 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U791 ( .A1(n703), .A2(n919), .ZN(n704) );
  XOR2_X1 U792 ( .A(KEYINPUT28), .B(n704), .Z(n705) );
  NOR2_X2 U793 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U794 ( .A(n707), .B(KEYINPUT29), .ZN(n713) );
  XNOR2_X1 U795 ( .A(G2078), .B(KEYINPUT93), .ZN(n708) );
  XNOR2_X1 U796 ( .A(n708), .B(KEYINPUT25), .ZN(n978) );
  NOR2_X1 U797 ( .A1(n978), .A2(n724), .ZN(n711) );
  NOR2_X1 U798 ( .A1(n709), .A2(G1961), .ZN(n710) );
  NOR2_X1 U799 ( .A1(n711), .A2(n710), .ZN(n718) );
  OR2_X1 U800 ( .A1(G301), .A2(n718), .ZN(n712) );
  NAND2_X1 U801 ( .A1(n713), .A2(n712), .ZN(n723) );
  NOR2_X1 U802 ( .A1(G1966), .A2(n797), .ZN(n737) );
  NOR2_X1 U803 ( .A1(G2084), .A2(n724), .ZN(n734) );
  NOR2_X1 U804 ( .A1(n737), .A2(n734), .ZN(n714) );
  NAND2_X1 U805 ( .A1(G8), .A2(n714), .ZN(n715) );
  XNOR2_X1 U806 ( .A(KEYINPUT30), .B(n715), .ZN(n716) );
  NOR2_X1 U807 ( .A1(G168), .A2(n716), .ZN(n717) );
  XNOR2_X1 U808 ( .A(n717), .B(KEYINPUT97), .ZN(n720) );
  NAND2_X1 U809 ( .A1(n718), .A2(G301), .ZN(n719) );
  NAND2_X1 U810 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U811 ( .A(n721), .B(KEYINPUT31), .ZN(n722) );
  NAND2_X1 U812 ( .A1(n723), .A2(n722), .ZN(n735) );
  NAND2_X1 U813 ( .A1(n735), .A2(G286), .ZN(n731) );
  INV_X1 U814 ( .A(G8), .ZN(n729) );
  NOR2_X1 U815 ( .A1(G1971), .A2(n797), .ZN(n726) );
  NOR2_X1 U816 ( .A1(G2090), .A2(n724), .ZN(n725) );
  NOR2_X1 U817 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U818 ( .A1(n727), .A2(G303), .ZN(n728) );
  OR2_X1 U819 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n733) );
  INV_X1 U821 ( .A(KEYINPUT32), .ZN(n732) );
  XNOR2_X1 U822 ( .A(n733), .B(n732), .ZN(n741) );
  NAND2_X1 U823 ( .A1(G8), .A2(n734), .ZN(n739) );
  INV_X1 U824 ( .A(n735), .ZN(n736) );
  NOR2_X1 U825 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U827 ( .A1(n741), .A2(n740), .ZN(n742) );
  XNOR2_X2 U828 ( .A(n742), .B(KEYINPUT98), .ZN(n763) );
  NOR2_X1 U829 ( .A1(G1971), .A2(G303), .ZN(n928) );
  NOR2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n743) );
  XOR2_X1 U831 ( .A(KEYINPUT99), .B(n743), .Z(n922) );
  NOR2_X1 U832 ( .A1(n928), .A2(n922), .ZN(n744) );
  NAND2_X1 U833 ( .A1(n763), .A2(n744), .ZN(n745) );
  XOR2_X1 U834 ( .A(KEYINPUT100), .B(n745), .Z(n746) );
  NOR2_X1 U835 ( .A1(n797), .A2(n746), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n925), .A2(n747), .ZN(n748) );
  NOR2_X1 U837 ( .A1(KEYINPUT101), .A2(n748), .ZN(n773) );
  NOR2_X1 U838 ( .A1(n750), .A2(n749), .ZN(n816) );
  XNOR2_X1 U839 ( .A(G2067), .B(KEYINPUT37), .ZN(n814) );
  XNOR2_X1 U840 ( .A(KEYINPUT86), .B(KEYINPUT34), .ZN(n754) );
  NAND2_X1 U841 ( .A1(n893), .A2(G140), .ZN(n752) );
  NAND2_X1 U842 ( .A1(G104), .A2(n666), .ZN(n751) );
  NAND2_X1 U843 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U844 ( .A(n754), .B(n753), .ZN(n760) );
  XNOR2_X1 U845 ( .A(KEYINPUT87), .B(KEYINPUT35), .ZN(n758) );
  NAND2_X1 U846 ( .A1(G128), .A2(n887), .ZN(n756) );
  NAND2_X1 U847 ( .A1(G116), .A2(n888), .ZN(n755) );
  NAND2_X1 U848 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U849 ( .A(n758), .B(n757), .ZN(n759) );
  NOR2_X1 U850 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U851 ( .A(n761), .B(KEYINPUT36), .ZN(n879) );
  NOR2_X1 U852 ( .A1(n814), .A2(n879), .ZN(n1005) );
  NAND2_X1 U853 ( .A1(n816), .A2(n1005), .ZN(n811) );
  NOR2_X1 U854 ( .A1(G2090), .A2(G303), .ZN(n762) );
  NAND2_X1 U855 ( .A1(G8), .A2(n762), .ZN(n764) );
  NAND2_X1 U856 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U857 ( .A1(n765), .A2(n797), .ZN(n770) );
  NOR2_X1 U858 ( .A1(G1981), .A2(G305), .ZN(n766) );
  XOR2_X1 U859 ( .A(n766), .B(KEYINPUT24), .Z(n767) );
  XNOR2_X1 U860 ( .A(KEYINPUT92), .B(n767), .ZN(n768) );
  OR2_X1 U861 ( .A1(n797), .A2(n768), .ZN(n769) );
  NAND2_X1 U862 ( .A1(n770), .A2(n769), .ZN(n771) );
  AND2_X1 U863 ( .A1(n811), .A2(n771), .ZN(n801) );
  OR2_X1 U864 ( .A1(KEYINPUT33), .A2(n801), .ZN(n772) );
  OR2_X1 U865 ( .A1(n773), .A2(n772), .ZN(n805) );
  XOR2_X1 U866 ( .A(G1986), .B(G290), .Z(n926) );
  XOR2_X1 U867 ( .A(KEYINPUT89), .B(G1991), .Z(n979) );
  NAND2_X1 U868 ( .A1(n893), .A2(G131), .ZN(n775) );
  NAND2_X1 U869 ( .A1(G95), .A2(n666), .ZN(n774) );
  NAND2_X1 U870 ( .A1(n775), .A2(n774), .ZN(n776) );
  XOR2_X1 U871 ( .A(KEYINPUT88), .B(n776), .Z(n780) );
  NAND2_X1 U872 ( .A1(G119), .A2(n887), .ZN(n778) );
  NAND2_X1 U873 ( .A1(G107), .A2(n888), .ZN(n777) );
  AND2_X1 U874 ( .A1(n778), .A2(n777), .ZN(n779) );
  NAND2_X1 U875 ( .A1(n780), .A2(n779), .ZN(n878) );
  NAND2_X1 U876 ( .A1(n979), .A2(n878), .ZN(n789) );
  NAND2_X1 U877 ( .A1(G129), .A2(n887), .ZN(n782) );
  NAND2_X1 U878 ( .A1(G117), .A2(n888), .ZN(n781) );
  NAND2_X1 U879 ( .A1(n782), .A2(n781), .ZN(n785) );
  NAND2_X1 U880 ( .A1(n666), .A2(G105), .ZN(n783) );
  XOR2_X1 U881 ( .A(KEYINPUT38), .B(n783), .Z(n784) );
  NOR2_X1 U882 ( .A1(n785), .A2(n784), .ZN(n787) );
  NAND2_X1 U883 ( .A1(n893), .A2(G141), .ZN(n786) );
  NAND2_X1 U884 ( .A1(n787), .A2(n786), .ZN(n884) );
  NAND2_X1 U885 ( .A1(G1996), .A2(n884), .ZN(n788) );
  NAND2_X1 U886 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U887 ( .A(KEYINPUT90), .B(n790), .Z(n806) );
  NAND2_X1 U888 ( .A1(n926), .A2(n806), .ZN(n791) );
  NAND2_X1 U889 ( .A1(n791), .A2(n816), .ZN(n803) );
  XOR2_X1 U890 ( .A(G1981), .B(G305), .Z(n936) );
  AND2_X1 U891 ( .A1(n936), .A2(n811), .ZN(n799) );
  INV_X1 U892 ( .A(KEYINPUT101), .ZN(n793) );
  NAND2_X1 U893 ( .A1(n922), .A2(KEYINPUT33), .ZN(n792) );
  NAND2_X1 U894 ( .A1(n793), .A2(n792), .ZN(n795) );
  NAND2_X1 U895 ( .A1(n922), .A2(KEYINPUT101), .ZN(n794) );
  NAND2_X1 U896 ( .A1(n795), .A2(n794), .ZN(n796) );
  OR2_X1 U897 ( .A1(n797), .A2(n796), .ZN(n798) );
  AND2_X1 U898 ( .A1(n799), .A2(n798), .ZN(n800) );
  OR2_X1 U899 ( .A1(n801), .A2(n800), .ZN(n802) );
  AND2_X1 U900 ( .A1(n803), .A2(n802), .ZN(n804) );
  NAND2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n819) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n884), .ZN(n1001) );
  INV_X1 U903 ( .A(n806), .ZN(n1009) );
  NOR2_X1 U904 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U905 ( .A1(n979), .A2(n878), .ZN(n997) );
  NOR2_X1 U906 ( .A1(n807), .A2(n997), .ZN(n808) );
  NOR2_X1 U907 ( .A1(n1009), .A2(n808), .ZN(n809) );
  NOR2_X1 U908 ( .A1(n1001), .A2(n809), .ZN(n810) );
  XNOR2_X1 U909 ( .A(n810), .B(KEYINPUT39), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U911 ( .A(n813), .B(KEYINPUT102), .ZN(n815) );
  NAND2_X1 U912 ( .A1(n814), .A2(n879), .ZN(n1011) );
  NAND2_X1 U913 ( .A1(n815), .A2(n1011), .ZN(n817) );
  NAND2_X1 U914 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U916 ( .A(KEYINPUT40), .B(n820), .ZN(G329) );
  XNOR2_X1 U917 ( .A(G2427), .B(G2435), .ZN(n830) );
  XOR2_X1 U918 ( .A(G2454), .B(G2430), .Z(n822) );
  XNOR2_X1 U919 ( .A(G2443), .B(G2451), .ZN(n821) );
  XNOR2_X1 U920 ( .A(n822), .B(n821), .ZN(n826) );
  XOR2_X1 U921 ( .A(G2446), .B(KEYINPUT103), .Z(n824) );
  XNOR2_X1 U922 ( .A(G1348), .B(G1341), .ZN(n823) );
  XNOR2_X1 U923 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U924 ( .A(n826), .B(n825), .Z(n828) );
  XNOR2_X1 U925 ( .A(G2438), .B(KEYINPUT104), .ZN(n827) );
  XNOR2_X1 U926 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U927 ( .A(n830), .B(n829), .ZN(n831) );
  NAND2_X1 U928 ( .A1(n831), .A2(G14), .ZN(n912) );
  XNOR2_X1 U929 ( .A(KEYINPUT105), .B(n912), .ZN(G401) );
  NAND2_X1 U930 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U931 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U932 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U933 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U934 ( .A1(n835), .A2(n834), .ZN(G188) );
  NAND2_X1 U936 ( .A1(n837), .A2(n836), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(G145) );
  INV_X1 U938 ( .A(G96), .ZN(G221) );
  INV_X1 U939 ( .A(G57), .ZN(G237) );
  NOR2_X1 U940 ( .A1(n841), .A2(n840), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U942 ( .A(G1956), .B(KEYINPUT41), .ZN(n851) );
  XOR2_X1 U943 ( .A(G1976), .B(G1981), .Z(n843) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1961), .ZN(n842) );
  XNOR2_X1 U945 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U946 ( .A(G1986), .B(G1991), .Z(n845) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1971), .ZN(n844) );
  XNOR2_X1 U948 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U949 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U950 ( .A(G2474), .B(KEYINPUT108), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(G229) );
  XOR2_X1 U953 ( .A(G2678), .B(KEYINPUT106), .Z(n853) );
  XNOR2_X1 U954 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n852) );
  XNOR2_X1 U955 ( .A(n853), .B(n852), .ZN(n857) );
  XOR2_X1 U956 ( .A(KEYINPUT42), .B(G2067), .Z(n855) );
  XNOR2_X1 U957 ( .A(G2090), .B(G2072), .ZN(n854) );
  XNOR2_X1 U958 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U959 ( .A(n857), .B(n856), .Z(n859) );
  XNOR2_X1 U960 ( .A(G2096), .B(G2100), .ZN(n858) );
  XNOR2_X1 U961 ( .A(n859), .B(n858), .ZN(n861) );
  XOR2_X1 U962 ( .A(G2078), .B(G2084), .Z(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(G227) );
  INV_X1 U964 ( .A(n862), .ZN(G319) );
  NAND2_X1 U965 ( .A1(n887), .A2(G124), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U967 ( .A1(G112), .A2(n888), .ZN(n864) );
  NAND2_X1 U968 ( .A1(n865), .A2(n864), .ZN(n869) );
  NAND2_X1 U969 ( .A1(n893), .A2(G136), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G100), .A2(n666), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n868) );
  NOR2_X1 U972 ( .A1(n869), .A2(n868), .ZN(G162) );
  NAND2_X1 U973 ( .A1(n893), .A2(G139), .ZN(n871) );
  NAND2_X1 U974 ( .A1(G103), .A2(n666), .ZN(n870) );
  NAND2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G127), .A2(n887), .ZN(n873) );
  NAND2_X1 U977 ( .A1(G115), .A2(n888), .ZN(n872) );
  NAND2_X1 U978 ( .A1(n873), .A2(n872), .ZN(n874) );
  XOR2_X1 U979 ( .A(KEYINPUT47), .B(n874), .Z(n875) );
  NOR2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n1013) );
  XOR2_X1 U981 ( .A(G164), .B(n1013), .Z(n877) );
  XNOR2_X1 U982 ( .A(n878), .B(n877), .ZN(n883) );
  XNOR2_X1 U983 ( .A(KEYINPUT48), .B(KEYINPUT111), .ZN(n881) );
  XNOR2_X1 U984 ( .A(n879), .B(KEYINPUT46), .ZN(n880) );
  XNOR2_X1 U985 ( .A(n881), .B(n880), .ZN(n882) );
  XNOR2_X1 U986 ( .A(n883), .B(n882), .ZN(n886) );
  XNOR2_X1 U987 ( .A(n884), .B(G162), .ZN(n885) );
  XNOR2_X1 U988 ( .A(n886), .B(n885), .ZN(n900) );
  NAND2_X1 U989 ( .A1(G130), .A2(n887), .ZN(n890) );
  NAND2_X1 U990 ( .A1(G118), .A2(n888), .ZN(n889) );
  NAND2_X1 U991 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U992 ( .A(KEYINPUT109), .B(n891), .Z(n898) );
  NAND2_X1 U993 ( .A1(G106), .A2(n666), .ZN(n892) );
  XNOR2_X1 U994 ( .A(n892), .B(KEYINPUT110), .ZN(n895) );
  NAND2_X1 U995 ( .A1(G142), .A2(n893), .ZN(n894) );
  NAND2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U997 ( .A(n896), .B(KEYINPUT45), .Z(n897) );
  NOR2_X1 U998 ( .A1(n898), .A2(n897), .ZN(n899) );
  XOR2_X1 U999 ( .A(n900), .B(n899), .Z(n902) );
  XNOR2_X1 U1000 ( .A(n994), .B(G160), .ZN(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n903), .ZN(G395) );
  XOR2_X1 U1003 ( .A(KEYINPUT112), .B(n904), .Z(n906) );
  XNOR2_X1 U1004 ( .A(G171), .B(G286), .ZN(n905) );
  XNOR2_X1 U1005 ( .A(n906), .B(n905), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n941), .B(n918), .ZN(n907) );
  XNOR2_X1 U1007 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n909), .ZN(G397) );
  NOR2_X1 U1009 ( .A1(G229), .A2(G227), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n910) );
  XNOR2_X1 U1011 ( .A(n911), .B(n910), .ZN(n915) );
  NAND2_X1 U1012 ( .A1(G319), .A2(n912), .ZN(n913) );
  XOR2_X1 U1013 ( .A(KEYINPUT113), .B(n913), .Z(n914) );
  NOR2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1018 ( .A(n918), .B(G1348), .Z(n934) );
  XOR2_X1 U1019 ( .A(G1956), .B(n919), .Z(n921) );
  NAND2_X1 U1020 ( .A1(G1971), .A2(G303), .ZN(n920) );
  NAND2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n932) );
  XNOR2_X1 U1022 ( .A(G301), .B(G1961), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(n922), .B(KEYINPUT124), .ZN(n923) );
  NOR2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n930) );
  NAND2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(KEYINPUT125), .B(n935), .ZN(n940) );
  XNOR2_X1 U1031 ( .A(G1966), .B(G168), .ZN(n937) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1033 ( .A(n938), .B(KEYINPUT57), .ZN(n939) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n943) );
  XNOR2_X1 U1035 ( .A(G1341), .B(n941), .ZN(n942) );
  NOR2_X1 U1036 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1037 ( .A(KEYINPUT126), .B(n944), .Z(n946) );
  XNOR2_X1 U1038 ( .A(G16), .B(KEYINPUT56), .ZN(n945) );
  NAND2_X1 U1039 ( .A1(n946), .A2(n945), .ZN(n1029) );
  XNOR2_X1 U1040 ( .A(G1348), .B(KEYINPUT59), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(n947), .B(G4), .ZN(n951) );
  XNOR2_X1 U1042 ( .A(G1956), .B(G20), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(G1341), .B(G19), .ZN(n948) );
  NOR2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n954) );
  XOR2_X1 U1046 ( .A(KEYINPUT127), .B(G1981), .Z(n952) );
  XNOR2_X1 U1047 ( .A(G6), .B(n952), .ZN(n953) );
  NOR2_X1 U1048 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(KEYINPUT60), .B(n955), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(G1966), .B(G21), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(G5), .B(G1961), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n966) );
  XNOR2_X1 U1054 ( .A(G1971), .B(G22), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(G23), .B(G1976), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n963) );
  XOR2_X1 U1057 ( .A(G1986), .B(G24), .Z(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(KEYINPUT58), .B(n964), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(KEYINPUT61), .B(n967), .ZN(n969) );
  INV_X1 U1062 ( .A(G16), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n970), .A2(G11), .ZN(n1027) );
  XOR2_X1 U1065 ( .A(G2090), .B(G35), .Z(n973) );
  XOR2_X1 U1066 ( .A(KEYINPUT54), .B(G34), .Z(n971) );
  XNOR2_X1 U1067 ( .A(n971), .B(G2084), .ZN(n972) );
  NAND2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n990) );
  XNOR2_X1 U1069 ( .A(G1996), .B(KEYINPUT121), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(n974), .B(G32), .ZN(n975) );
  NAND2_X1 U1071 ( .A1(n975), .A2(G28), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(G33), .B(G2072), .ZN(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n983) );
  XNOR2_X1 U1074 ( .A(n978), .B(G27), .ZN(n981) );
  XNOR2_X1 U1075 ( .A(n979), .B(G25), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(KEYINPUT120), .B(G2067), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(G26), .B(n984), .ZN(n985) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1081 ( .A(KEYINPUT53), .B(n987), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(KEYINPUT122), .B(n988), .ZN(n989) );
  NOR2_X1 U1083 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1084 ( .A(KEYINPUT55), .B(n991), .Z(n992) );
  NOR2_X1 U1085 ( .A1(G29), .A2(n992), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(n993), .B(KEYINPUT123), .ZN(n1025) );
  XNOR2_X1 U1087 ( .A(G160), .B(G2084), .ZN(n995) );
  NAND2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n1007) );
  XNOR2_X1 U1090 ( .A(KEYINPUT117), .B(KEYINPUT51), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(n998), .B(KEYINPUT116), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G2090), .B(G162), .ZN(n999) );
  XNOR2_X1 U1093 ( .A(n999), .B(KEYINPUT115), .ZN(n1000) );
  NOR2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1095 ( .A(n1003), .B(n1002), .Z(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(n1010), .B(KEYINPUT118), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XNOR2_X1 U1101 ( .A(G2072), .B(n1013), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(G164), .B(G2078), .ZN(n1014) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1104 ( .A(KEYINPUT119), .B(n1016), .Z(n1017) );
  XNOR2_X1 U1105 ( .A(KEYINPUT50), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1107 ( .A(n1020), .B(KEYINPUT52), .ZN(n1022) );
  INV_X1 U1108 ( .A(KEYINPUT55), .ZN(n1021) );
  NAND2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(G29), .A2(n1023), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1030), .Z(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

