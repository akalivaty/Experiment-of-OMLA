//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:38 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n557, new_n558,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1191, new_n1192;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT64), .ZN(G220));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XOR2_X1   g014(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XOR2_X1   g019(.A(new_n444), .B(KEYINPUT67), .Z(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G219), .A4(G221), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n463), .A2(G137), .A3(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n466), .A2(G2105), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  AND2_X1   g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n470), .B1(new_n463), .B2(G125), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT68), .B1(new_n471), .B2(new_n464), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  NOR2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n473), .B(G2105), .C1(new_n478), .C2(new_n470), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n469), .B1(new_n472), .B2(new_n479), .ZN(G160));
  INV_X1    g055(.A(new_n463), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n481), .A2(new_n464), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n464), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  AND2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  OAI211_X1 g065(.A(G138), .B(new_n464), .C1(new_n490), .C2(new_n475), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n463), .A2(new_n493), .A3(G138), .A4(new_n464), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OR2_X1    g070(.A1(G102), .A2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(G2105), .B1(KEYINPUT69), .B2(G114), .ZN(new_n497));
  AND2_X1   g072(.A1(KEYINPUT69), .A2(G114), .ZN(new_n498));
  OAI211_X1 g073(.A(G2104), .B(new_n496), .C1(new_n497), .C2(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G126), .B(G2105), .C1(new_n490), .C2(new_n475), .ZN(new_n500));
  AND2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  AND2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT6), .A2(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n506), .A2(G88), .B1(G50), .B2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n504), .A2(G62), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(new_n511), .B1(KEYINPUT70), .B2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(new_n515), .A2(KEYINPUT70), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n516), .A2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  INV_X1    g095(.A(G51), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n505), .A2(G543), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  AND2_X1   g098(.A1(G63), .A2(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n504), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n523), .B1(new_n504), .B2(new_n524), .ZN(new_n527));
  OAI221_X1 g102(.A(new_n520), .B1(new_n521), .B2(new_n522), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n529), .A2(KEYINPUT73), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(KEYINPUT73), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(KEYINPUT7), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT7), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n530), .A2(new_n534), .A3(new_n531), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n533), .A2(new_n535), .B1(G89), .B2(new_n506), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n526), .A2(new_n527), .B1(new_n521), .B2(new_n522), .ZN(new_n538));
  AND2_X1   g113(.A1(new_n538), .A2(KEYINPUT72), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n537), .A2(new_n539), .ZN(G168));
  AOI22_X1  g115(.A1(new_n506), .A2(G90), .B1(G52), .B2(new_n510), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n504), .A2(G64), .ZN(new_n542));
  NAND2_X1  g117(.A1(G77), .A2(G543), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n512), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n541), .B1(KEYINPUT74), .B2(new_n544), .ZN(new_n545));
  AND2_X1   g120(.A1(new_n544), .A2(KEYINPUT74), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n545), .A2(new_n546), .ZN(G171));
  NAND2_X1  g122(.A1(new_n504), .A2(new_n505), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n548), .A2(new_n549), .B1(new_n522), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n512), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(new_n510), .A2(G53), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n548), .A2(KEYINPUT75), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT75), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n504), .A2(new_n505), .A3(new_n563), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(G91), .A3(new_n564), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n566));
  OR2_X1    g141(.A1(new_n566), .A2(new_n512), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n561), .A2(new_n565), .A3(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  NAND3_X1  g145(.A1(new_n562), .A2(G87), .A3(new_n564), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n504), .A2(G74), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G651), .B1(G49), .B2(new_n510), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(G288));
  NAND2_X1  g149(.A1(new_n504), .A2(G61), .ZN(new_n575));
  NAND2_X1  g150(.A1(G73), .A2(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(G48), .B2(new_n510), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n562), .A2(G86), .A3(new_n564), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(G305));
  INV_X1    g155(.A(G85), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n548), .A2(new_n581), .B1(new_n522), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n584), .A2(new_n512), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G290));
  NAND2_X1  g162(.A1(G301), .A2(G868), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n562), .A2(G92), .A3(new_n564), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(KEYINPUT76), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n591));
  NAND4_X1  g166(.A1(new_n562), .A2(new_n591), .A3(G92), .A4(new_n564), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n590), .A2(KEYINPUT10), .A3(new_n592), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n504), .A2(G66), .ZN(new_n597));
  INV_X1    g172(.A(G79), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n507), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n599), .A2(G651), .B1(G54), .B2(new_n510), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n595), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n588), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n588), .B1(new_n602), .B2(G868), .ZN(G321));
  INV_X1    g179(.A(G868), .ZN(new_n605));
  NOR2_X1   g180(.A1(G168), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  AND3_X1   g182(.A1(new_n561), .A2(new_n565), .A3(new_n567), .ZN(new_n608));
  OAI211_X1 g183(.A(new_n607), .B(KEYINPUT77), .C1(G868), .C2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(KEYINPUT77), .B2(new_n607), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT78), .ZN(G297));
  XNOR2_X1  g186(.A(new_n610), .B(KEYINPUT79), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n602), .B1(new_n613), .B2(G860), .ZN(G148));
  INV_X1    g189(.A(new_n554), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(new_n605), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n601), .A2(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(new_n605), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g194(.A1(new_n463), .A2(new_n467), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT12), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT13), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G2100), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT80), .Z(new_n624));
  NAND2_X1  g199(.A1(new_n482), .A2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n484), .A2(G123), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n464), .A2(G111), .ZN(new_n627));
  OAI21_X1  g202(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT81), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2096), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n624), .B(new_n631), .C1(G2100), .C2(new_n622), .ZN(G156));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2427), .B(G2430), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n636), .A2(KEYINPUT14), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT82), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(new_n634), .B2(new_n635), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n643), .A2(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n646), .A2(new_n647), .A3(G14), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G401));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2072), .B(G2078), .Z(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT18), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n653), .B(KEYINPUT17), .ZN(new_n656));
  INV_X1    g231(.A(new_n650), .ZN(new_n657));
  INV_X1    g232(.A(new_n651), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n656), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n653), .A3(new_n658), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(new_n652), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n655), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT20), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n667), .A2(new_n668), .ZN(new_n672));
  NOR3_X1   g247(.A1(new_n666), .A2(new_n669), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n673), .B1(new_n666), .B2(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(G1981), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT83), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n679), .A2(new_n681), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  OR3_X1    g260(.A1(new_n682), .A2(new_n683), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n682), .B2(new_n683), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(G229));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n689), .A2(G25), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(KEYINPUT84), .Z(new_n691));
  AOI22_X1  g266(.A1(G119), .A2(new_n484), .B1(new_n482), .B2(G131), .ZN(new_n692));
  INV_X1    g267(.A(G95), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(new_n464), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT85), .ZN(new_n695));
  OAI21_X1  g270(.A(G2104), .B1(new_n464), .B2(G107), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n692), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT86), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n691), .B1(new_n698), .B2(G29), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT87), .Z(new_n700));
  XOR2_X1   g275(.A(KEYINPUT35), .B(G1991), .Z(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  AND2_X1   g277(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n700), .A2(new_n702), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT88), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(KEYINPUT88), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n708), .A2(G24), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n586), .B(KEYINPUT89), .Z(new_n710));
  AOI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n708), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1986), .ZN(new_n712));
  NOR3_X1   g287(.A1(new_n703), .A2(new_n704), .A3(new_n712), .ZN(new_n713));
  MUX2_X1   g288(.A(G6), .B(G305), .S(G16), .Z(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT90), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT32), .B(G1981), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n708), .ZN(new_n718));
  NOR2_X1   g293(.A1(G166), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G22), .B2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G1971), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  MUX2_X1   g298(.A(G23), .B(G288), .S(G16), .Z(new_n724));
  XOR2_X1   g299(.A(KEYINPUT33), .B(G1976), .Z(new_n725));
  XOR2_X1   g300(.A(new_n724), .B(new_n725), .Z(new_n726));
  NAND4_X1  g301(.A1(new_n717), .A2(new_n722), .A3(new_n723), .A4(new_n726), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n727), .A2(KEYINPUT34), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n713), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT91), .B(KEYINPUT36), .Z(new_n731));
  OR2_X1    g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n689), .A2(G32), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n484), .A2(G129), .ZN(new_n735));
  NAND3_X1  g310(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT26), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n482), .A2(G141), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n467), .A2(G105), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n734), .B1(new_n742), .B2(new_n689), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT27), .B(G1996), .Z(new_n744));
  NOR2_X1   g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g320(.A1(new_n689), .A2(G33), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n482), .A2(G139), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT93), .ZN(new_n748));
  NAND3_X1  g323(.A1(new_n464), .A2(G103), .A3(G2104), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT25), .Z(new_n750));
  AOI22_X1  g325(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n748), .B(new_n750), .C1(new_n464), .C2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n746), .B1(new_n752), .B2(G29), .ZN(new_n753));
  INV_X1    g328(.A(G2072), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n745), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g330(.A(new_n755), .B1(new_n754), .B2(new_n753), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT24), .ZN(new_n757));
  INV_X1    g332(.A(G34), .ZN(new_n758));
  AOI21_X1  g333(.A(G29), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n757), .B2(new_n758), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G160), .B2(new_n689), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n756), .B1(G2084), .B2(new_n761), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT94), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n718), .A2(G20), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT23), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n608), .B2(new_n705), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT98), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1956), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n602), .A2(G16), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G4), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT92), .B(G1348), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n768), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G29), .A2(G35), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G162), .B2(G29), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT97), .B(KEYINPUT29), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2090), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n689), .A2(G26), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT28), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n482), .A2(G140), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n484), .A2(G128), .ZN(new_n781));
  OR2_X1    g356(.A1(G104), .A2(G2105), .ZN(new_n782));
  OAI211_X1 g357(.A(new_n782), .B(G2104), .C1(G116), .C2(new_n464), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n779), .B1(new_n785), .B2(new_n689), .ZN(new_n786));
  INV_X1    g361(.A(G2067), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  XOR2_X1   g363(.A(KEYINPUT31), .B(G11), .Z(new_n789));
  INV_X1    g364(.A(KEYINPUT30), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n689), .B1(new_n790), .B2(G28), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT95), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n791), .A2(new_n792), .B1(new_n790), .B2(G28), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n789), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n629), .B2(new_n689), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n743), .B2(new_n744), .ZN(new_n797));
  OAI211_X1 g372(.A(new_n788), .B(new_n797), .C1(G2084), .C2(new_n761), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n777), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n689), .A2(G27), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G164), .B2(new_n689), .ZN(new_n801));
  INV_X1    g376(.A(G2078), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n708), .A2(G19), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(new_n554), .B2(new_n708), .ZN(new_n805));
  INV_X1    g380(.A(G1341), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n803), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n705), .A2(G5), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G171), .B2(new_n705), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1961), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n705), .A2(G21), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G168), .B2(new_n705), .ZN(new_n813));
  AOI211_X1 g388(.A(new_n808), .B(new_n811), .C1(G1966), .C2(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(G1966), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT96), .Z(new_n816));
  NAND2_X1  g391(.A1(new_n770), .A2(new_n771), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n799), .A2(new_n814), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n763), .A2(new_n772), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n732), .A2(new_n733), .A3(new_n819), .ZN(G150));
  INV_X1    g395(.A(G150), .ZN(G311));
  NAND2_X1  g396(.A1(new_n602), .A2(G559), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT38), .ZN(new_n823));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  INV_X1    g399(.A(G55), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n548), .A2(new_n824), .B1(new_n522), .B2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT99), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(new_n512), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n827), .A2(new_n554), .A3(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n554), .B1(new_n827), .B2(new_n829), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n823), .B(new_n833), .ZN(new_n834));
  AND2_X1   g409(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n834), .A2(KEYINPUT39), .ZN(new_n836));
  NOR3_X1   g411(.A1(new_n835), .A2(new_n836), .A3(G860), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n827), .A2(new_n829), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(G860), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n837), .A2(new_n840), .ZN(G145));
  XNOR2_X1  g416(.A(G162), .B(new_n629), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(G160), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n499), .A2(new_n500), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n844), .A2(KEYINPUT100), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT100), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n499), .A2(new_n500), .A3(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n495), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n784), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n752), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n742), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n697), .B(new_n621), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n482), .A2(G142), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n484), .A2(G130), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT101), .ZN(new_n856));
  INV_X1    g431(.A(G118), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n855), .A2(new_n856), .B1(new_n857), .B2(G2105), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n856), .B2(new_n855), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n853), .A2(new_n854), .A3(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n852), .B(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(new_n851), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(KEYINPUT102), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n851), .A2(new_n861), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n862), .A2(KEYINPUT102), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n843), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(KEYINPUT103), .B(G37), .Z(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n843), .B1(new_n851), .B2(new_n861), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n869), .B1(new_n862), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g448(.A1(new_n838), .A2(new_n605), .ZN(new_n874));
  XOR2_X1   g449(.A(G303), .B(G305), .Z(new_n875));
  XNOR2_X1  g450(.A(G288), .B(new_n586), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n875), .B(new_n876), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT42), .ZN(new_n878));
  OR2_X1    g453(.A1(new_n831), .A2(new_n832), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n617), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n596), .A2(new_n600), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT10), .B1(new_n590), .B2(new_n592), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n608), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND4_X1  g458(.A1(new_n595), .A2(G299), .A3(new_n596), .A4(new_n600), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT104), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n883), .A2(new_n888), .A3(new_n884), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT41), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n601), .A2(KEYINPUT104), .A3(new_n608), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n883), .A2(KEYINPUT41), .A3(new_n884), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT106), .A4(KEYINPUT41), .ZN(new_n896));
  AOI22_X1  g471(.A1(new_n892), .A2(KEYINPUT105), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT105), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n889), .A2(new_n898), .A3(new_n890), .A4(new_n891), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n887), .B1(new_n900), .B2(new_n880), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n878), .B(new_n901), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n874), .B1(new_n902), .B2(new_n605), .ZN(G295));
  OAI21_X1  g478(.A(new_n874), .B1(new_n902), .B2(new_n605), .ZN(G331));
  INV_X1    g479(.A(KEYINPUT110), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT107), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n537), .B2(new_n539), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n538), .A2(KEYINPUT72), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n908), .A2(KEYINPUT107), .A3(new_n528), .A4(new_n536), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n907), .A2(G301), .A3(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(G168), .A2(KEYINPUT107), .A3(G171), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n879), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n833), .A2(new_n911), .A3(new_n910), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n890), .B1(new_n889), .B2(new_n891), .ZN(new_n916));
  OAI22_X1  g491(.A1(new_n916), .A2(KEYINPUT109), .B1(KEYINPUT41), .B2(new_n886), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT109), .ZN(new_n918));
  AOI211_X1 g493(.A(new_n918), .B(new_n890), .C1(new_n889), .C2(new_n891), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n915), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n913), .A2(new_n914), .A3(new_n921), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n833), .A2(KEYINPUT108), .A3(new_n911), .A4(new_n910), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n885), .ZN(new_n925));
  AND2_X1   g500(.A1(new_n920), .A2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n877), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n905), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT43), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n927), .B1(new_n920), .B2(new_n925), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT110), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n915), .A2(new_n886), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n922), .A2(new_n923), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n932), .B1(new_n900), .B2(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n869), .B1(new_n934), .B2(new_n927), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n928), .A2(new_n929), .A3(new_n931), .A4(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(G37), .B1(new_n934), .B2(new_n927), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n924), .B1(new_n899), .B2(new_n897), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n877), .B1(new_n938), .B2(new_n932), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT44), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n900), .A2(new_n933), .ZN(new_n945));
  INV_X1    g520(.A(new_n932), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n945), .A2(new_n927), .A3(new_n946), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n947), .B(new_n868), .C1(new_n930), .C2(KEYINPUT110), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n930), .A2(KEYINPUT110), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT43), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G37), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n939), .A2(new_n947), .A3(new_n929), .A4(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT111), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n937), .A2(KEYINPUT111), .A3(new_n929), .A4(new_n939), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n950), .A2(KEYINPUT44), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n944), .A2(new_n956), .ZN(G397));
  INV_X1    g532(.A(KEYINPUT123), .ZN(new_n958));
  INV_X1    g533(.A(G1384), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n848), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT45), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G40), .ZN(new_n963));
  AOI211_X1 g538(.A(new_n963), .B(new_n469), .C1(new_n472), .C2(new_n479), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n502), .A2(new_n959), .ZN(new_n965));
  OAI211_X1 g540(.A(new_n962), .B(new_n964), .C1(new_n961), .C2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(G1966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(KEYINPUT50), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT50), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n848), .A2(new_n970), .A3(new_n959), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n964), .A3(new_n971), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n972), .A2(G2084), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n968), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(G8), .B1(new_n974), .B2(G286), .ZN(new_n975));
  AND2_X1   g550(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(KEYINPUT122), .A2(KEYINPUT51), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  OAI211_X1 g554(.A(G8), .B(new_n979), .C1(new_n974), .C2(G286), .ZN(new_n980));
  INV_X1    g555(.A(G8), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(new_n968), .B2(new_n973), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(G286), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n977), .A2(new_n980), .A3(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT117), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n970), .B1(new_n848), .B2(new_n959), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n472), .A2(new_n479), .ZN(new_n987));
  INV_X1    g562(.A(new_n469), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n987), .A2(G40), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n985), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  AOI22_X1  g565(.A1(KEYINPUT100), .A2(new_n844), .B1(new_n492), .B2(new_n494), .ZN(new_n991));
  AOI21_X1  g566(.A(G1384), .B1(new_n991), .B2(new_n847), .ZN(new_n992));
  OAI211_X1 g567(.A(new_n964), .B(KEYINPUT117), .C1(new_n992), .C2(new_n970), .ZN(new_n993));
  INV_X1    g568(.A(G2090), .ZN(new_n994));
  AOI21_X1  g569(.A(G1384), .B1(new_n495), .B2(new_n501), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n970), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n990), .A2(new_n993), .A3(new_n994), .A4(new_n996), .ZN(new_n997));
  XOR2_X1   g572(.A(KEYINPUT113), .B(G1971), .Z(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n965), .A2(new_n961), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n964), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n960), .A2(new_n961), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n999), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n981), .B1(new_n997), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(G303), .A2(G8), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT55), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n964), .A2(new_n992), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n571), .A2(new_n573), .A3(G1976), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(G8), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(KEYINPUT52), .ZN(new_n1014));
  INV_X1    g589(.A(G1976), .ZN(new_n1015));
  AOI21_X1  g590(.A(KEYINPUT52), .B1(G288), .B2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1011), .A2(G8), .A3(new_n1016), .A4(new_n1012), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n578), .A2(new_n579), .A3(new_n676), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(KEYINPUT115), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n578), .A2(new_n579), .A3(new_n1021), .A4(new_n676), .ZN(new_n1022));
  INV_X1    g597(.A(G86), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n578), .B1(new_n1023), .B2(new_n548), .ZN(new_n1024));
  AOI22_X1  g599(.A1(new_n1020), .A2(new_n1022), .B1(G1981), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT49), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1011), .A2(G8), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1024), .A2(G1981), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT49), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n1027), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1018), .B1(new_n1026), .B2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n995), .A2(KEYINPUT45), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1034), .A2(new_n989), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n992), .A2(KEYINPUT45), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n998), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n969), .A2(new_n971), .A3(new_n964), .A4(new_n994), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT114), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT114), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1003), .A2(new_n1041), .A3(new_n1038), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1040), .A2(new_n1042), .A3(new_n1009), .A4(G8), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1033), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1035), .A2(new_n802), .A3(new_n1036), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n1046));
  INV_X1    g621(.A(G1961), .ZN(new_n1047));
  AOI22_X1  g622(.A1(new_n1045), .A2(new_n1046), .B1(new_n1047), .B2(new_n972), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1046), .A2(G2078), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n966), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g627(.A(G171), .B(KEYINPUT54), .Z(new_n1053));
  INV_X1    g628(.A(new_n962), .ZN(new_n1054));
  NOR3_X1   g629(.A1(new_n469), .A2(new_n963), .A3(new_n1050), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n464), .B2(new_n471), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1054), .A2(new_n1002), .A3(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1053), .A2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n1052), .A2(new_n1053), .B1(new_n1058), .B2(new_n1048), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n984), .A2(new_n1010), .A3(new_n1044), .A4(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(new_n608), .B(KEYINPUT57), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1063));
  XOR2_X1   g638(.A(KEYINPUT56), .B(G2072), .Z(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n990), .A2(new_n993), .A3(new_n996), .ZN(new_n1067));
  INV_X1    g642(.A(G1956), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(KEYINPUT119), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(KEYINPUT119), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1066), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT119), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1065), .B1(new_n1075), .B2(new_n1069), .ZN(new_n1076));
  OAI211_X1 g651(.A(KEYINPUT61), .B(new_n1072), .C1(new_n1076), .C2(new_n1061), .ZN(new_n1077));
  INV_X1    g652(.A(G1996), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1036), .A2(new_n1078), .A3(new_n964), .A4(new_n1000), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1080));
  XNOR2_X1  g655(.A(new_n1080), .B(new_n806), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1011), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n615), .B1(new_n1079), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1084), .A2(KEYINPUT121), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1083), .B(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G1348), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n972), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n989), .A2(new_n960), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(new_n787), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(new_n602), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n601), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT60), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OR3_X1    g670(.A1(new_n1092), .A2(KEYINPUT60), .A3(new_n601), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1087), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1098), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1075), .A2(new_n1069), .ZN(new_n1100));
  AOI22_X1  g675(.A1(new_n1099), .A2(new_n1062), .B1(new_n1100), .B2(new_n1066), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1077), .B(new_n1097), .C1(new_n1101), .C2(KEYINPUT61), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1076), .A2(new_n1061), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1072), .B1(new_n1103), .B2(new_n1094), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1060), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT118), .B(KEYINPUT63), .Z(new_n1106));
  OAI211_X1 g681(.A(new_n1033), .B(new_n1043), .C1(new_n1009), .C2(new_n1004), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n982), .A2(G168), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1108), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1040), .A2(G8), .A3(new_n1042), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1111), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1044), .A2(KEYINPUT63), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1109), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n571), .A2(new_n573), .A3(new_n1015), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n1032), .B2(new_n1026), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1028), .ZN(new_n1117));
  OAI21_X1  g692(.A(KEYINPUT116), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT116), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1090), .A2(new_n981), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n1025), .B2(KEYINPUT49), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  OAI211_X1 g698(.A(new_n1119), .B(new_n1028), .C1(new_n1123), .C2(new_n1115), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1118), .A2(new_n1124), .A3(new_n1120), .ZN(new_n1125));
  OR3_X1    g700(.A1(new_n1043), .A2(new_n1123), .A3(new_n1018), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1114), .A2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n958), .B1(new_n1105), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1098), .A2(new_n1061), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(new_n1075), .B2(new_n1069), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1099), .A2(new_n1062), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1094), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1087), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT61), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1133), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1139), .B2(new_n1134), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1138), .B1(new_n1103), .B2(new_n1133), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1136), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n1131), .B(KEYINPUT123), .C1(new_n1142), .C2(new_n1060), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1044), .A2(G171), .A3(new_n1010), .A4(new_n1052), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT124), .ZN(new_n1146));
  OAI211_X1 g721(.A(new_n1145), .B(new_n1146), .C1(KEYINPUT62), .C2(new_n984), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n984), .A2(KEYINPUT62), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT124), .B1(new_n1148), .B2(new_n1144), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n984), .A2(KEYINPUT62), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1147), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1129), .A2(new_n1143), .A3(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n962), .A2(new_n989), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n1078), .ZN(new_n1154));
  XNOR2_X1  g729(.A(new_n1154), .B(KEYINPUT112), .ZN(new_n1155));
  INV_X1    g730(.A(new_n742), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1153), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n784), .B(new_n787), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1156), .A2(G1996), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n697), .B(new_n701), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1162), .B1(new_n1158), .B2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n586), .B(new_n678), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1164), .B1(new_n1153), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1152), .A2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n784), .A2(G2067), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n698), .A2(new_n702), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1168), .B1(new_n1162), .B2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NOR4_X1   g747(.A1(new_n1157), .A2(new_n698), .A3(new_n702), .A4(new_n1161), .ZN(new_n1173));
  OAI21_X1  g748(.A(KEYINPUT125), .B1(new_n1173), .B2(new_n1168), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1172), .A2(new_n1174), .A3(KEYINPUT126), .A4(new_n1153), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1172), .A2(new_n1174), .A3(new_n1153), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT126), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n1159), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1153), .B1(new_n1179), .B2(new_n1156), .ZN(new_n1180));
  AND2_X1   g755(.A1(new_n1155), .A2(KEYINPUT46), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n1155), .A2(KEYINPUT46), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g758(.A(new_n1183), .B(KEYINPUT47), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1153), .A2(new_n678), .A3(new_n586), .ZN(new_n1185));
  XOR2_X1   g760(.A(new_n1185), .B(KEYINPUT48), .Z(new_n1186));
  OR2_X1    g761(.A1(new_n1164), .A2(new_n1186), .ZN(new_n1187));
  AND4_X1   g762(.A1(new_n1175), .A2(new_n1178), .A3(new_n1184), .A4(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1167), .A2(new_n1188), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g764(.A1(new_n461), .A2(G227), .ZN(new_n1191));
  NOR3_X1   g765(.A1(G229), .A2(G401), .A3(new_n1191), .ZN(new_n1192));
  AND3_X1   g766(.A1(new_n942), .A2(new_n1192), .A3(new_n872), .ZN(G308));
  NAND3_X1  g767(.A1(new_n942), .A2(new_n1192), .A3(new_n872), .ZN(G225));
endmodule


