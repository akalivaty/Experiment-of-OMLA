//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 1 0 1 0 1 0 0 0 1 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1273, new_n1274, new_n1275,
    new_n1276;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n210), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(new_n201), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n227));
  INV_X1    g0027(.A(G58), .ZN(new_n228));
  INV_X1    g0028(.A(G232), .ZN(new_n229));
  INV_X1    g0029(.A(G257), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n205), .C2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n212), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n215), .B1(new_n218), .B2(new_n220), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(new_n229), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G58), .B(G77), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT64), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XOR2_X1   g0047(.A(G107), .B(G116), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n216), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(new_n202), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n210), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(G77), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n256), .A2(new_n257), .B1(new_n210), .B2(G68), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n252), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT11), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n252), .B1(new_n209), .B2(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G68), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT12), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n264), .B1(new_n266), .B2(new_n222), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n265), .A2(KEYINPUT12), .A3(G68), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n263), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n259), .A2(new_n260), .ZN(new_n270));
  NOR3_X1   g0070(.A1(new_n261), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G274), .ZN(new_n275));
  INV_X1    g0075(.A(G33), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  OAI211_X1 g0077(.A(G1), .B(G13), .C1(new_n276), .C2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(new_n273), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n275), .B1(new_n279), .B2(new_n223), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT67), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n280), .B(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n287), .A2(G232), .B1(G33), .B2(G97), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT3), .B(G33), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(G226), .A3(new_n286), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XOR2_X1   g0093(.A(KEYINPUT68), .B(KEYINPUT13), .Z(new_n294));
  NAND3_X1  g0094(.A1(new_n282), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n280), .B(KEYINPUT67), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n278), .B1(new_n288), .B2(new_n290), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT13), .ZN(new_n299));
  OAI211_X1 g0099(.A(new_n295), .B(G179), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G169), .ZN(new_n301));
  INV_X1    g0101(.A(new_n294), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(new_n296), .B2(new_n297), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(new_n303), .B2(new_n295), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT14), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n300), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AOI211_X1 g0106(.A(KEYINPUT14), .B(new_n301), .C1(new_n303), .C2(new_n295), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n272), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n295), .B(G190), .C1(new_n298), .C2(new_n299), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n303), .A2(new_n295), .ZN(new_n310));
  INV_X1    g0110(.A(G200), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n271), .B(new_n309), .C1(new_n310), .C2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT3), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n276), .ZN(new_n316));
  NAND2_X1  g0116(.A1(KEYINPUT3), .A2(G33), .ZN(new_n317));
  AOI21_X1  g0117(.A(G1698), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G222), .ZN(new_n319));
  INV_X1    g0119(.A(G223), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n289), .A2(G1698), .ZN(new_n321));
  OAI221_X1 g0121(.A(new_n319), .B1(new_n257), .B2(new_n289), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n292), .ZN(new_n323));
  INV_X1    g0123(.A(new_n275), .ZN(new_n324));
  INV_X1    g0124(.A(new_n279), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n324), .B1(new_n325), .B2(G226), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n323), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(G200), .ZN(new_n328));
  XOR2_X1   g0128(.A(new_n328), .B(KEYINPUT66), .Z(new_n329));
  INV_X1    g0129(.A(new_n252), .ZN(new_n330));
  XNOR2_X1  g0130(.A(KEYINPUT8), .B(G58), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT65), .ZN(new_n332));
  XNOR2_X1  g0132(.A(new_n331), .B(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n256), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n253), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n330), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n262), .A2(G50), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n338), .B1(G50), .B2(new_n265), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  OR2_X1    g0140(.A1(new_n340), .A2(KEYINPUT9), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(KEYINPUT9), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n323), .A2(G190), .A3(new_n326), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT10), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n329), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  XNOR2_X1  g0146(.A(new_n328), .B(KEYINPUT66), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT10), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n340), .B1(new_n301), .B2(new_n327), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n323), .A2(new_n352), .A3(new_n326), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n325), .A2(G244), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n318), .A2(G232), .ZN(new_n357));
  OAI221_X1 g0157(.A(new_n357), .B1(new_n206), .B2(new_n289), .C1(new_n223), .C2(new_n321), .ZN(new_n358));
  AOI211_X1 g0158(.A(new_n324), .B(new_n356), .C1(new_n358), .C2(new_n292), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n359), .A2(new_n352), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n262), .A2(G77), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT15), .B(G87), .ZN(new_n362));
  INV_X1    g0162(.A(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n363), .A2(new_n334), .B1(G20), .B2(G77), .ZN(new_n364));
  OR2_X1    g0164(.A1(new_n331), .A2(new_n254), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI221_X1 g0166(.A(new_n361), .B1(G77), .B2(new_n265), .C1(new_n366), .C2(new_n330), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n359), .B2(G169), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n367), .B1(new_n359), .B2(G190), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n311), .B2(new_n359), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n314), .A2(new_n350), .A3(new_n355), .A4(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(G223), .B(new_n286), .C1(new_n283), .C2(new_n284), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT71), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n289), .A2(KEYINPUT71), .A3(G223), .A4(new_n286), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  OAI211_X1 g0179(.A(G226), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n380));
  NAND2_X1  g0180(.A1(G33), .A2(G87), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n278), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n275), .B1(new_n279), .B2(new_n229), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n311), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G190), .ZN(new_n387));
  INV_X1    g0187(.A(new_n385), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n382), .B1(new_n377), .B2(new_n378), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n387), .B(new_n388), .C1(new_n389), .C2(new_n278), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT73), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NOR2_X1   g0193(.A1(new_n228), .A2(new_n222), .ZN(new_n394));
  OAI21_X1  g0194(.A(G20), .B1(new_n394), .B2(new_n201), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n253), .A2(G159), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n316), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n317), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT69), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(new_n283), .B2(new_n284), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n316), .A2(KEYINPUT69), .A3(new_n317), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n402), .A2(new_n403), .A3(new_n210), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n400), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(KEYINPUT16), .B(new_n398), .C1(new_n406), .C2(new_n222), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT70), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n399), .A2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n285), .A2(KEYINPUT70), .A3(KEYINPUT7), .A4(new_n210), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n405), .B1(new_n289), .B2(G20), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n397), .B1(new_n412), .B2(G68), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n407), .B(new_n252), .C1(new_n413), .C2(KEYINPUT16), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n333), .A2(new_n265), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n333), .B2(new_n262), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n386), .A2(KEYINPUT73), .A3(new_n390), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n393), .A2(new_n414), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  XNOR2_X1  g0218(.A(new_n418), .B(KEYINPUT17), .ZN(new_n419));
  OAI21_X1  g0219(.A(G169), .B1(new_n384), .B2(new_n385), .ZN(new_n420));
  OAI211_X1 g0220(.A(G179), .B(new_n388), .C1(new_n389), .C2(new_n278), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT72), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n407), .A2(new_n252), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n413), .A2(KEYINPUT16), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n416), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n420), .A2(KEYINPUT72), .A3(new_n421), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n424), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT18), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n429), .B(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n419), .A2(new_n431), .ZN(new_n432));
  OR3_X1    g0232(.A1(new_n374), .A2(KEYINPUT74), .A3(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT74), .B1(new_n374), .B2(new_n432), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n318), .A2(KEYINPUT77), .A3(G250), .ZN(new_n436));
  OAI211_X1 g0236(.A(G250), .B(new_n286), .C1(new_n283), .C2(new_n284), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT77), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n289), .A2(G257), .A3(G1698), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G294), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n436), .A2(new_n439), .A3(new_n440), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n292), .ZN(new_n443));
  XNOR2_X1  g0243(.A(KEYINPUT5), .B(G41), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n209), .A2(G45), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n444), .A2(new_n278), .A3(G274), .A4(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n292), .B1(new_n446), .B2(new_n444), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G264), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n443), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G200), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n210), .B(G87), .C1(new_n283), .C2(new_n284), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(KEYINPUT22), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT22), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n289), .A2(new_n454), .A3(new_n210), .A4(G87), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G116), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n457), .A2(G20), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT23), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(new_n210), .B2(G107), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT24), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n330), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(new_n464), .B2(new_n463), .ZN(new_n466));
  OR3_X1    g0266(.A1(new_n265), .A2(KEYINPUT25), .A3(G107), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT25), .B1(new_n265), .B2(G107), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n209), .A2(G33), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n265), .A2(new_n469), .A3(new_n216), .A4(new_n251), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n467), .B(new_n468), .C1(new_n206), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT76), .ZN(new_n472));
  INV_X1    g0272(.A(new_n470), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G107), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT76), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n474), .A2(new_n475), .A3(new_n467), .A4(new_n468), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n442), .A2(new_n292), .B1(G264), .B2(new_n448), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n478), .A2(G190), .A3(new_n447), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n451), .A2(new_n466), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n460), .A2(new_n461), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n481), .B1(G20), .B2(new_n457), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(new_n453), .B2(new_n455), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n252), .B1(new_n483), .B2(KEYINPUT24), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n463), .A2(new_n464), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n477), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n450), .A2(new_n301), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n478), .A2(new_n352), .A3(new_n447), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n486), .A2(new_n487), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n480), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT78), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n480), .A2(new_n489), .A3(KEYINPUT78), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n266), .A2(new_n205), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(new_n470), .B2(new_n205), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n412), .A2(G107), .ZN(new_n497));
  XNOR2_X1  g0297(.A(G97), .B(G107), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT6), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n499), .A2(new_n205), .A3(G107), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n503), .A2(G20), .B1(G77), .B2(new_n253), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n497), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n496), .B1(new_n505), .B2(new_n252), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n444), .A2(new_n446), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n278), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n447), .B1(new_n508), .B2(new_n230), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n289), .A2(G244), .A3(new_n286), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT4), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(G33), .A2(G283), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n318), .A2(KEYINPUT4), .A3(G244), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n289), .A2(G250), .A3(G1698), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n512), .A2(new_n513), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n509), .B1(new_n516), .B2(new_n292), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G190), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n506), .B(new_n518), .C1(new_n311), .C2(new_n517), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n516), .A2(new_n292), .ZN(new_n520));
  INV_X1    g0320(.A(new_n509), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n301), .ZN(new_n523));
  INV_X1    g0323(.A(new_n496), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n501), .B1(new_n499), .B2(new_n498), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n525), .A2(new_n210), .B1(new_n257), .B2(new_n254), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n526), .B1(G107), .B2(new_n412), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n524), .B1(new_n527), .B2(new_n330), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n517), .A2(new_n352), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n523), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n445), .A2(G250), .ZN(new_n531));
  INV_X1    g0331(.A(G274), .ZN(new_n532));
  OAI22_X1  g0332(.A1(new_n292), .A2(new_n531), .B1(new_n532), .B2(new_n445), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n289), .A2(G238), .A3(new_n286), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n289), .A2(G244), .A3(G1698), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n534), .A2(new_n535), .A3(new_n457), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n533), .B1(new_n536), .B2(new_n292), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n289), .A2(new_n210), .A3(G68), .ZN(new_n538));
  NAND3_X1  g0338(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n210), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(G87), .B2(new_n207), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT19), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n542), .B1(new_n256), .B2(new_n205), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n538), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  AOI22_X1  g0344(.A1(new_n544), .A2(new_n252), .B1(new_n266), .B2(new_n362), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n473), .A2(new_n363), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n352), .A2(new_n537), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(new_n537), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n301), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  OR3_X1    g0350(.A1(new_n470), .A2(KEYINPUT75), .A3(new_n224), .ZN(new_n551));
  OAI21_X1  g0351(.A(KEYINPUT75), .B1(new_n470), .B2(new_n224), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n545), .A2(new_n553), .ZN(new_n554));
  AOI211_X1 g0354(.A(new_n387), .B(new_n533), .C1(new_n536), .C2(new_n292), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n548), .A2(G200), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n519), .A2(new_n530), .A3(new_n550), .A4(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(new_n513), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n560), .B(new_n252), .C1(new_n210), .C2(G116), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT20), .ZN(new_n562));
  XNOR2_X1  g0362(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(G116), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n266), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n473), .A2(G116), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n444), .A2(new_n446), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n292), .A2(new_n532), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n448), .A2(G270), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n289), .A2(G264), .A3(G1698), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n285), .A2(G303), .ZN(new_n573));
  OAI211_X1 g0373(.A(G257), .B(new_n286), .C1(new_n283), .C2(new_n284), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n292), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(G200), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n568), .B(new_n578), .C1(new_n387), .C2(new_n577), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT21), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(G169), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n568), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n567), .A2(KEYINPUT21), .A3(G169), .A4(new_n577), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n571), .A2(new_n576), .A3(G179), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n567), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n579), .A2(new_n582), .A3(new_n583), .A4(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n559), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n435), .A2(new_n494), .A3(new_n587), .ZN(G372));
  INV_X1    g0388(.A(KEYINPUT83), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n536), .A2(new_n292), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(KEYINPUT79), .ZN(new_n591));
  XNOR2_X1  g0391(.A(new_n533), .B(KEYINPUT80), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT79), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n536), .A2(new_n593), .A3(new_n292), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n547), .B1(new_n595), .B2(G169), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n556), .B1(new_n595), .B2(new_n311), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(new_n530), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n599), .A2(KEYINPUT26), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n558), .A2(new_n550), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n530), .ZN(new_n602));
  XNOR2_X1  g0402(.A(KEYINPUT82), .B(KEYINPUT26), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n589), .B(new_n596), .C1(new_n600), .C2(new_n604), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n523), .A2(new_n529), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(new_n596), .A3(new_n597), .A4(new_n528), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT26), .ZN(new_n608));
  AOI22_X1  g0408(.A1(new_n607), .A2(new_n608), .B1(new_n602), .B2(new_n603), .ZN(new_n609));
  INV_X1    g0409(.A(new_n596), .ZN(new_n610));
  OAI21_X1  g0410(.A(KEYINPUT83), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n480), .A2(new_n519), .A3(new_n530), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n612), .A2(new_n598), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT81), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT81), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n612), .B2(new_n598), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n582), .A2(new_n585), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n617), .A2(new_n489), .A3(new_n583), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n614), .A2(new_n616), .A3(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n605), .A2(new_n611), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n435), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n427), .A2(new_n422), .ZN(new_n622));
  XNOR2_X1  g0422(.A(new_n622), .B(new_n430), .ZN(new_n623));
  INV_X1    g0423(.A(new_n308), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n312), .B2(new_n369), .ZN(new_n625));
  INV_X1    g0425(.A(new_n419), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n354), .B1(new_n627), .B2(new_n350), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n621), .A2(new_n628), .ZN(G369));
  NAND3_X1  g0429(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n630));
  OR2_X1    g0430(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(KEYINPUT27), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n631), .A2(G213), .A3(new_n632), .ZN(new_n633));
  INV_X1    g0433(.A(G343), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n567), .A2(new_n635), .ZN(new_n636));
  XOR2_X1   g0436(.A(new_n636), .B(KEYINPUT84), .Z(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n617), .A2(new_n583), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n640), .B1(new_n586), .B2(new_n638), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(G330), .ZN(new_n642));
  INV_X1    g0442(.A(new_n635), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n489), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n486), .A2(new_n635), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n494), .B2(new_n645), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n639), .A2(new_n643), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n492), .B2(new_n493), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n635), .B(KEYINPUT85), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n489), .A2(new_n651), .ZN(new_n652));
  NOR2_X1   g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n648), .A2(new_n653), .ZN(G399));
  INV_X1    g0454(.A(new_n213), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n655), .A2(G41), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n224), .A2(new_n205), .A3(new_n206), .A4(new_n564), .ZN(new_n658));
  XOR2_X1   g0458(.A(new_n658), .B(KEYINPUT86), .Z(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n657), .A2(G1), .A3(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n661), .B1(new_n220), .B2(new_n657), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n662), .B(KEYINPUT28), .ZN(new_n663));
  INV_X1    g0463(.A(new_n651), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n494), .A2(new_n587), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT31), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n584), .A2(new_n517), .A3(new_n478), .A4(new_n537), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT87), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT30), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n443), .A2(new_n537), .A3(new_n449), .ZN(new_n671));
  NAND4_X1  g0471(.A1(new_n671), .A2(KEYINPUT30), .A3(new_n584), .A4(new_n517), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n591), .A2(new_n592), .A3(new_n594), .ZN(new_n673));
  AOI21_X1  g0473(.A(G179), .B1(new_n571), .B2(new_n576), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n673), .A2(new_n522), .A3(new_n450), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n668), .B1(new_n667), .B2(new_n669), .ZN(new_n677));
  NOR3_X1   g0477(.A1(new_n670), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n666), .B1(new_n678), .B2(new_n643), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n667), .A2(new_n669), .ZN(new_n680));
  OAI211_X1 g0480(.A(KEYINPUT31), .B(new_n651), .C1(new_n676), .C2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n665), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(G330), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n620), .A2(new_n664), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT88), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT29), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n620), .A2(KEYINPUT88), .A3(new_n664), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n687), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n602), .A2(new_n603), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n599), .A2(KEYINPUT26), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n610), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n613), .A2(new_n618), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n635), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(KEYINPUT29), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n684), .B1(new_n690), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n663), .B1(new_n697), .B2(G1), .ZN(G364));
  AND2_X1   g0498(.A1(new_n210), .A2(G13), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n209), .B1(new_n699), .B2(G45), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n656), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n216), .B1(G20), .B2(new_n301), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n210), .A2(new_n387), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n311), .A2(G179), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n352), .A2(G200), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  AOI22_X1  g0512(.A1(G303), .A2(new_n709), .B1(new_n712), .B2(G322), .ZN(new_n713));
  INV_X1    g0513(.A(G311), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n210), .A2(G190), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n710), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n713), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n352), .A2(new_n311), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n706), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(KEYINPUT91), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n719), .A2(KEYINPUT91), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n717), .B1(G326), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(G179), .A2(G200), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G190), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G20), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G294), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n718), .A2(new_n715), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  XNOR2_X1  g0531(.A(KEYINPUT33), .B(G317), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n289), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n715), .A2(new_n707), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n715), .A2(new_n726), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI22_X1  g0537(.A1(G283), .A2(new_n735), .B1(new_n737), .B2(G329), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n725), .A2(new_n729), .A3(new_n733), .A4(new_n738), .ZN(new_n739));
  XOR2_X1   g0539(.A(new_n739), .B(KEYINPUT92), .Z(new_n740));
  NOR2_X1   g0540(.A1(new_n708), .A2(new_n224), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(G107), .B2(new_n735), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n742), .B(new_n289), .C1(new_n222), .C2(new_n730), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n743), .B1(G50), .B2(new_n724), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n728), .A2(G97), .ZN(new_n745));
  INV_X1    g0545(.A(G159), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n736), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT32), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n711), .A2(new_n228), .B1(new_n716), .B2(new_n257), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT90), .ZN(new_n750));
  NAND4_X1  g0550(.A1(new_n744), .A2(new_n745), .A3(new_n748), .A4(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(new_n705), .B1(new_n740), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(G13), .A2(G33), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n704), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n213), .A2(new_n289), .ZN(new_n757));
  INV_X1    g0557(.A(G355), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n757), .A2(new_n758), .B1(G116), .B2(new_n213), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT89), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n245), .A2(G45), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n402), .A2(new_n403), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n655), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(G45), .B2(new_n220), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n760), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n703), .B(new_n752), .C1(new_n756), .C2(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(new_n755), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n766), .B1(new_n641), .B2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n641), .A2(G330), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n642), .A2(new_n703), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT93), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(G396));
  NAND2_X1  g0573(.A1(new_n367), .A2(new_n635), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n372), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(new_n370), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n369), .A2(new_n643), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n687), .A2(new_n689), .A3(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n778), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n620), .A2(new_n664), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g0581(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n684), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n782), .A2(new_n684), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n784), .A2(new_n703), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n783), .B1(new_n785), .B2(KEYINPUT97), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(KEYINPUT97), .B2(new_n785), .ZN(new_n787));
  INV_X1    g0587(.A(new_n716), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G143), .A2(new_n712), .B1(new_n788), .B2(G159), .ZN(new_n789));
  INV_X1    g0589(.A(G150), .ZN(new_n790));
  INV_X1    g0590(.A(G137), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n789), .B1(new_n790), .B2(new_n730), .C1(new_n723), .C2(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(KEYINPUT94), .B(KEYINPUT34), .Z(new_n793));
  XNOR2_X1  g0593(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n735), .A2(G68), .ZN(new_n795));
  INV_X1    g0595(.A(new_n728), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n795), .B1(new_n202), .B2(new_n708), .C1(new_n228), .C2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n762), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(G132), .B2(new_n737), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n797), .B1(new_n799), .B2(KEYINPUT95), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n794), .B(new_n800), .C1(KEYINPUT95), .C2(new_n799), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n724), .A2(G303), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n716), .A2(new_n564), .B1(new_n736), .B2(new_n714), .ZN(new_n803));
  AOI211_X1 g0603(.A(new_n289), .B(new_n803), .C1(G87), .C2(new_n735), .ZN(new_n804));
  INV_X1    g0604(.A(G294), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n206), .A2(new_n708), .B1(new_n711), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G283), .B2(new_n731), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n802), .A2(new_n804), .A3(new_n745), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n705), .B1(new_n801), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n704), .A2(new_n753), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n703), .B(new_n809), .C1(new_n257), .C2(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(new_n811), .B(KEYINPUT96), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n754), .B2(new_n780), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n787), .A2(new_n813), .ZN(G384));
  AOI211_X1 g0614(.A(new_n564), .B(new_n218), .C1(new_n503), .C2(KEYINPUT35), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(KEYINPUT35), .B2(new_n503), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT36), .Z(new_n817));
  OR3_X1    g0617(.A1(new_n220), .A2(new_n257), .A3(new_n394), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n202), .A2(G68), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n209), .B(G13), .C1(new_n818), .C2(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT39), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT38), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT17), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n418), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(new_n417), .ZN(new_n826));
  AOI21_X1  g0626(.A(KEYINPUT73), .B1(new_n386), .B2(new_n390), .ZN(new_n827));
  NOR3_X1   g0627(.A1(new_n826), .A2(new_n427), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(KEYINPUT17), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n623), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  AOI211_X1 g0630(.A(KEYINPUT100), .B(new_n633), .C1(new_n414), .C2(new_n416), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT100), .ZN(new_n832));
  INV_X1    g0632(.A(new_n633), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n427), .B2(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n830), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT99), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n424), .A2(new_n427), .A3(new_n837), .A4(new_n428), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  AND3_X1   g0640(.A1(new_n420), .A2(KEYINPUT72), .A3(new_n421), .ZN(new_n841));
  AOI21_X1  g0641(.A(KEYINPUT72), .B1(new_n420), .B2(new_n421), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n837), .B1(new_n843), .B2(new_n427), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n831), .ZN(new_n846));
  INV_X1    g0646(.A(new_n834), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n828), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n418), .B(new_n622), .C1(new_n831), .C2(new_n834), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n845), .A2(new_n848), .B1(KEYINPUT37), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n836), .B1(new_n850), .B2(KEYINPUT101), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n849), .A2(KEYINPUT37), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n418), .B1(new_n831), .B2(new_n834), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n853), .A2(new_n844), .A3(new_n840), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT101), .ZN(new_n855));
  NOR3_X1   g0655(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  OAI211_X1 g0656(.A(KEYINPUT102), .B(new_n823), .C1(new_n851), .C2(new_n856), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n406), .A2(new_n222), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT16), .B1(new_n858), .B2(new_n398), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n416), .B1(new_n859), .B2(new_n425), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n833), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n419), .B2(new_n431), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n861), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n860), .A2(new_n422), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n418), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n864), .B1(new_n866), .B2(KEYINPUT98), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT98), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n418), .A2(new_n865), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n839), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n863), .B(KEYINPUT38), .C1(new_n854), .C2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n857), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n850), .A2(KEYINPUT101), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n855), .B1(new_n852), .B2(new_n854), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n873), .A2(new_n874), .A3(new_n836), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT102), .B1(new_n875), .B2(new_n823), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n822), .B1(new_n872), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n870), .A2(new_n854), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n823), .B1(new_n878), .B2(new_n862), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(new_n871), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(new_n822), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n624), .A2(new_n643), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n877), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(new_n623), .A2(new_n833), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n271), .A2(new_n643), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n306), .B2(new_n307), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n313), .B2(new_n887), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n781), .B2(new_n777), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n886), .B1(new_n891), .B2(new_n880), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n885), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n690), .A2(new_n435), .A3(new_n696), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n628), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n893), .B(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(G330), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n676), .A2(new_n677), .ZN(new_n898));
  OAI211_X1 g0698(.A(KEYINPUT31), .B(new_n635), .C1(new_n898), .C2(new_n670), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n665), .A2(new_n679), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(new_n889), .A3(new_n780), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(KEYINPUT40), .B1(new_n880), .B2(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n823), .B1(new_n851), .B2(new_n856), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT102), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n906), .A2(new_n857), .A3(new_n871), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n901), .A2(KEYINPUT103), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT103), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n900), .A2(new_n889), .A3(new_n780), .A4(new_n909), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n908), .A2(KEYINPUT40), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n903), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n435), .A2(new_n900), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n897), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n915), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n896), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n209), .B2(new_n699), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n896), .A2(new_n916), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n821), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT104), .ZN(G367));
  OAI211_X1 g0721(.A(new_n519), .B(new_n530), .C1(new_n506), .C2(new_n664), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n606), .A2(new_n528), .A3(new_n651), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n650), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n530), .B1(new_n922), .B2(new_n489), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n925), .A2(KEYINPUT42), .B1(new_n664), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n927), .B(KEYINPUT105), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n925), .A2(KEYINPUT42), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(KEYINPUT106), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n643), .B1(new_n545), .B2(new_n553), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n610), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n598), .B2(new_n932), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n930), .A2(KEYINPUT106), .A3(new_n934), .ZN(new_n937));
  NAND4_X1  g0737(.A1(new_n936), .A2(KEYINPUT43), .A3(new_n930), .A4(new_n937), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n936), .A2(new_n937), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n938), .B1(new_n939), .B2(KEYINPUT43), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n647), .A2(new_n924), .ZN(new_n941));
  OR2_X1    g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n656), .B(KEYINPUT41), .Z(new_n944));
  INV_X1    g0744(.A(new_n650), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n646), .A2(new_n649), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n945), .A2(new_n946), .A3(KEYINPUT107), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(KEYINPUT107), .B2(new_n946), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(new_n642), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n697), .A2(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n950), .A2(KEYINPUT108), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n653), .A2(new_n924), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT45), .Z(new_n953));
  NOR2_X1   g0753(.A1(new_n653), .A2(new_n924), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT44), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(new_n648), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n950), .A2(KEYINPUT108), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n951), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n944), .B1(new_n959), .B2(new_n697), .ZN(new_n960));
  OAI211_X1 g0760(.A(new_n942), .B(new_n943), .C1(new_n701), .C2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n763), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n756), .B1(new_n213), .B2(new_n362), .C1(new_n962), .C2(new_n241), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n963), .A2(new_n702), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT46), .ZN(new_n965));
  NOR3_X1   g0765(.A1(new_n708), .A2(new_n965), .A3(new_n564), .ZN(new_n966));
  INV_X1    g0766(.A(G303), .ZN(new_n967));
  INV_X1    g0767(.A(G317), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n798), .B1(new_n967), .B2(new_n711), .C1(new_n968), .C2(new_n736), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n966), .B(new_n969), .C1(G107), .C2(new_n728), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n965), .B1(new_n708), .B2(new_n564), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT109), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n735), .A2(G97), .ZN(new_n973));
  INV_X1    g0773(.A(G283), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n973), .B1(new_n974), .B2(new_n716), .C1(new_n805), .C2(new_n730), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G311), .B2(new_n724), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n970), .A2(new_n972), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n724), .A2(G143), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n730), .A2(new_n746), .B1(new_n736), .B2(new_n791), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n285), .B(new_n979), .C1(G58), .C2(new_n709), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n796), .A2(new_n222), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n711), .A2(new_n790), .B1(new_n716), .B2(new_n202), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n734), .A2(new_n257), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n978), .A2(new_n980), .A3(new_n982), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n977), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT47), .Z(new_n988));
  OAI221_X1 g0788(.A(new_n964), .B1(new_n934), .B2(new_n767), .C1(new_n988), .C2(new_n705), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n961), .A2(new_n989), .ZN(G387));
  NAND2_X1  g0790(.A1(new_n646), .A2(new_n755), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n660), .A2(new_n757), .B1(G107), .B2(new_n213), .ZN(new_n992));
  AOI211_X1 g0792(.A(G45), .B(new_n659), .C1(G68), .C2(G77), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(KEYINPUT110), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(KEYINPUT110), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n331), .A2(G50), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT50), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n994), .A2(new_n995), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n962), .B1(new_n238), .B2(G45), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n992), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(new_n756), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n702), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G311), .A2(new_n731), .B1(new_n788), .B2(G303), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n968), .B2(new_n711), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1004), .B1(G322), .B2(new_n724), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT48), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(KEYINPUT48), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n709), .A2(G294), .B1(new_n728), .B2(G283), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT49), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n734), .A2(new_n564), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n762), .B(new_n1012), .C1(G326), .C2(new_n737), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n796), .A2(new_n362), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n788), .A2(G68), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1016), .A2(new_n762), .A3(new_n973), .A4(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n708), .A2(new_n257), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(G50), .B2(new_n712), .ZN(new_n1020));
  XOR2_X1   g0820(.A(KEYINPUT111), .B(G150), .Z(new_n1021));
  OAI21_X1  g0821(.A(new_n1020), .B1(new_n736), .B2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(G159), .B2(new_n724), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n333), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1023), .B1(new_n1024), .B2(new_n730), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1011), .A2(new_n1014), .B1(new_n1018), .B2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1002), .B1(new_n1026), .B2(new_n704), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n949), .A2(new_n701), .B1(new_n991), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n950), .A2(new_n656), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n697), .A2(new_n949), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(G393));
  INV_X1    g0831(.A(new_n950), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n959), .B(new_n656), .C1(new_n1032), .C2(new_n957), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n957), .A2(new_n701), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n756), .B1(new_n205), .B2(new_n213), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1035), .B1(new_n763), .B2(new_n249), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n703), .A2(new_n1036), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n723), .A2(new_n790), .B1(new_n746), .B2(new_n711), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT51), .Z(new_n1039));
  AOI22_X1  g0839(.A1(G68), .A2(new_n709), .B1(new_n735), .B2(G87), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n737), .A2(G143), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1040), .A2(new_n762), .A3(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT112), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n796), .A2(new_n257), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n730), .A2(new_n202), .B1(new_n716), .B2(new_n331), .ZN(new_n1045));
  NOR4_X1   g0845(.A1(new_n1039), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n723), .A2(new_n968), .B1(new_n714), .B2(new_n711), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT52), .Z(new_n1048));
  AOI22_X1  g0848(.A1(G283), .A2(new_n709), .B1(new_n737), .B2(G322), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n805), .B2(new_n716), .C1(new_n967), .C2(new_n730), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n285), .B1(new_n734), .B2(new_n206), .C1(new_n796), .C2(new_n564), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n1048), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n1046), .A2(new_n1052), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1037), .B1(new_n767), .B2(new_n924), .C1(new_n1053), .C2(new_n705), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1033), .A2(new_n1034), .A3(new_n1054), .ZN(G390));
  NAND3_X1  g0855(.A1(new_n900), .A2(G330), .A3(new_n780), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1056), .A2(new_n890), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n891), .A2(new_n884), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n877), .B2(new_n882), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n695), .A2(new_n776), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n777), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n884), .B1(new_n1062), .B2(new_n889), .ZN(new_n1063));
  AND2_X1   g0863(.A1(new_n907), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1058), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n683), .A2(new_n778), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(new_n889), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n907), .A2(new_n1063), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n881), .B1(new_n907), .B2(new_n822), .ZN(new_n1069));
  OAI211_X1 g0869(.A(new_n1067), .B(new_n1068), .C1(new_n1069), .C2(new_n1059), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n1065), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n701), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n810), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n702), .B1(new_n333), .B2(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n795), .B1(new_n564), .B2(new_n711), .C1(new_n805), .C2(new_n736), .ZN(new_n1075));
  NOR4_X1   g0875(.A1(new_n1075), .A2(new_n289), .A3(new_n741), .A4(new_n1044), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G107), .A2(new_n731), .B1(new_n788), .B2(G97), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1077), .A2(KEYINPUT117), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n724), .A2(G283), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1077), .A2(KEYINPUT117), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1076), .A2(new_n1078), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1021), .A2(new_n708), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT53), .Z(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G159), .B2(new_n728), .ZN(new_n1084));
  INV_X1    g0884(.A(G125), .ZN(new_n1085));
  OAI221_X1 g0885(.A(new_n289), .B1(new_n736), .B2(new_n1085), .C1(new_n202), .C2(new_n734), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT115), .ZN(new_n1087));
  XNOR2_X1  g0887(.A(KEYINPUT54), .B(G143), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n730), .A2(new_n791), .B1(new_n716), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1086), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1084), .B(new_n1090), .C1(new_n1087), .C2(new_n1089), .ZN(new_n1091));
  INV_X1    g0891(.A(G128), .ZN(new_n1092));
  INV_X1    g0892(.A(G132), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n723), .A2(new_n1092), .B1(new_n1093), .B2(new_n711), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT116), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1081), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  OR2_X1    g0896(.A1(new_n1096), .A2(KEYINPUT118), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n705), .B1(new_n1096), .B2(KEYINPUT118), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1074), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n1069), .B2(new_n754), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1072), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n435), .A2(G330), .A3(new_n900), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n894), .A2(new_n628), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1056), .A2(new_n890), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1062), .B1(new_n889), .B2(new_n1066), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1057), .B1(new_n889), .B2(new_n1066), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n781), .A2(new_n777), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1105), .A2(new_n1106), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1065), .A2(new_n1070), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT113), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1065), .A2(new_n1070), .A3(new_n1110), .A4(KEYINPUT113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(KEYINPUT114), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1115), .A2(new_n1116), .A3(new_n656), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1071), .A2(new_n1110), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n657), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1121), .A2(new_n1116), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1102), .B1(new_n1120), .B2(new_n1122), .ZN(G378));
  OAI21_X1  g0923(.A(new_n702), .B1(G50), .B2(new_n1073), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n798), .A2(new_n277), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n724), .B2(G116), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1019), .B(new_n981), .C1(G107), .C2(new_n712), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n730), .A2(new_n205), .B1(new_n734), .B2(new_n228), .ZN(new_n1128));
  OAI22_X1  g0928(.A1(new_n716), .A2(new_n362), .B1(new_n736), .B2(new_n974), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1126), .A2(new_n1127), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT58), .ZN(new_n1132));
  AOI21_X1  g0932(.A(G50), .B1(new_n276), .B2(new_n277), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1131), .A2(new_n1132), .B1(new_n1125), .B2(new_n1133), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n730), .A2(new_n1093), .B1(new_n716), .B2(new_n791), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1092), .A2(new_n711), .B1(new_n708), .B2(new_n1088), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n1135), .B(new_n1136), .C1(G150), .C2(new_n728), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n1085), .B2(new_n723), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(KEYINPUT59), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n735), .A2(G159), .ZN(new_n1140));
  AOI211_X1 g0940(.A(G33), .B(G41), .C1(new_n737), .C2(G124), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1138), .A2(KEYINPUT59), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n1134), .B1(new_n1132), .B2(new_n1131), .C1(new_n1142), .C2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1124), .B1(new_n1144), .B2(new_n704), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n350), .A2(new_n355), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n340), .A2(new_n633), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1147), .B(KEYINPUT55), .ZN(new_n1148));
  XOR2_X1   g0948(.A(new_n1146), .B(new_n1148), .Z(new_n1149));
  XOR2_X1   g0949(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1150));
  XNOR2_X1  g0950(.A(new_n1149), .B(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1145), .B1(new_n1151), .B2(new_n754), .ZN(new_n1152));
  XOR2_X1   g0952(.A(new_n1152), .B(KEYINPUT120), .Z(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1151), .B1(new_n912), .B2(G330), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n911), .B1(new_n872), .B2(new_n876), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n880), .A2(new_n902), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT40), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AND4_X1   g0959(.A1(G330), .A2(new_n1156), .A3(new_n1151), .A4(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n893), .B1(new_n1155), .B2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1156), .A2(G330), .A3(new_n1159), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1151), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1156), .A2(new_n1151), .A3(G330), .A4(new_n1159), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1164), .A2(new_n885), .A3(new_n892), .A4(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT121), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1161), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(KEYINPUT121), .B(new_n893), .C1(new_n1155), .C2(new_n1160), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1154), .B1(new_n1170), .B2(new_n700), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1104), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1115), .A2(new_n1173), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1175));
  AOI21_X1  g0975(.A(KEYINPUT57), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1104), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1177));
  INV_X1    g0977(.A(KEYINPUT122), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1161), .A2(new_n1166), .A3(new_n1178), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n893), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1180), .A2(KEYINPUT122), .A3(new_n1165), .A4(new_n1164), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1179), .A2(KEYINPUT57), .A3(new_n1181), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n656), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1172), .B1(new_n1176), .B2(new_n1183), .ZN(G375));
  AOI21_X1  g0984(.A(new_n703), .B1(new_n222), .B2(new_n810), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT123), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n730), .A2(new_n564), .B1(new_n716), .B2(new_n206), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n723), .A2(new_n805), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(G97), .A2(new_n709), .B1(new_n712), .B2(G283), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1190), .B1(new_n967), .B2(new_n736), .ZN(new_n1191));
  NOR4_X1   g0991(.A1(new_n1191), .A2(new_n289), .A3(new_n984), .A4(new_n1015), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n711), .A2(new_n791), .B1(new_n736), .B2(new_n1092), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n746), .A2(new_n708), .B1(new_n730), .B2(new_n1088), .ZN(new_n1194));
  AOI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(new_n724), .C2(G132), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n228), .A2(new_n734), .B1(new_n716), .B2(new_n790), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n798), .B(new_n1196), .C1(G50), .C2(new_n728), .ZN(new_n1197));
  AOI22_X1  g0997(.A1(new_n1189), .A2(new_n1192), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n1185), .B1(new_n705), .B2(new_n1198), .C1(new_n889), .C2(new_n754), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1199), .B1(new_n1109), .B2(new_n700), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1104), .A2(new_n1109), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n944), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1201), .B1(new_n1203), .B2(new_n1205), .ZN(G381));
  AND3_X1   g1006(.A1(new_n1179), .A2(KEYINPUT57), .A3(new_n1181), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n657), .B1(new_n1174), .B2(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT57), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1177), .B2(new_n1170), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1171), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1121), .A2(new_n1116), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1118), .B1(new_n1121), .B2(new_n1116), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1101), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(G390), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n961), .A2(new_n989), .A3(new_n1216), .ZN(new_n1217));
  OR3_X1    g1017(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1218));
  OR4_X1    g1018(.A1(G381), .A2(new_n1215), .A3(new_n1217), .A4(new_n1218), .ZN(G407));
  OAI211_X1 g1019(.A(G407), .B(G213), .C1(G343), .C2(new_n1215), .ZN(G409));
  INV_X1    g1020(.A(KEYINPUT126), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(G393), .B(new_n772), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1217), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1216), .B1(new_n961), .B2(new_n989), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1221), .B(new_n1222), .C1(new_n1223), .C2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1224), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1222), .A2(new_n1221), .ZN(new_n1227));
  OR2_X1    g1027(.A1(new_n1222), .A2(new_n1221), .ZN(new_n1228));
  NAND4_X1  g1028(.A1(new_n1226), .A2(new_n1217), .A3(new_n1227), .A4(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1225), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT61), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n787), .A2(KEYINPUT125), .A3(new_n813), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT60), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1202), .B1(new_n1110), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1104), .A2(KEYINPUT60), .A3(new_n1109), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1234), .A2(new_n656), .A3(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1232), .A2(new_n1201), .A3(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT125), .B1(new_n787), .B2(new_n813), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT125), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1237), .A2(new_n1240), .A3(G384), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(G213), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(G343), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1244), .A2(G2897), .ZN(new_n1245));
  XNOR2_X1  g1045(.A(new_n1242), .B(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1179), .A2(new_n701), .A3(new_n1181), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1152), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1177), .A2(new_n1170), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1248), .B1(new_n1249), .B2(new_n1204), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(G378), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT124), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1252), .B1(G375), .B2(new_n1214), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1211), .A2(KEYINPUT124), .A3(G378), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1251), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1246), .B1(new_n1255), .B2(new_n1244), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1242), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1255), .A2(new_n1244), .A3(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT62), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1231), .B(new_n1256), .C1(new_n1258), .C2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1261));
  OR2_X1    g1061(.A1(G378), .A2(new_n1250), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1244), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1263), .A2(new_n1264), .A3(new_n1242), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1265), .A2(KEYINPUT62), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1230), .B1(new_n1260), .B2(new_n1266), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1230), .B1(new_n1258), .B2(KEYINPUT63), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT63), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1265), .A2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1268), .A2(new_n1231), .A3(new_n1270), .A4(new_n1256), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1267), .A2(new_n1271), .ZN(G405));
  NAND2_X1  g1072(.A1(G375), .A2(new_n1214), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1261), .A2(new_n1273), .ZN(new_n1274));
  XNOR2_X1  g1074(.A(new_n1274), .B(KEYINPUT127), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1230), .B(new_n1242), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1275), .B(new_n1276), .ZN(G402));
endmodule


