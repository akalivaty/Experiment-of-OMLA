//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n768, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G227), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n189), .B(KEYINPUT74), .ZN(new_n190));
  XNOR2_X1  g004(.A(G110), .B(G140), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT11), .ZN(new_n194));
  INV_X1    g008(.A(G134), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G137), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(KEYINPUT11), .A3(G134), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n195), .A2(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT66), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n202), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n204), .A2(new_n196), .A3(new_n198), .A4(new_n199), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT65), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  AND2_X1   g022(.A1(KEYINPUT64), .A2(G143), .ZN(new_n209));
  NOR2_X1   g023(.A1(KEYINPUT64), .A2(G143), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT1), .B1(new_n212), .B2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G128), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n212), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT64), .A2(G143), .ZN(new_n217));
  AOI21_X1  g031(.A(G146), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT65), .B1(new_n208), .B2(G143), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n211), .B(new_n214), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n212), .A2(G146), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G128), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n216), .A2(new_n217), .ZN(new_n225));
  OAI211_X1 g039(.A(new_n222), .B(new_n224), .C1(new_n225), .C2(new_n208), .ZN(new_n226));
  INV_X1    g040(.A(G107), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n227), .A2(G104), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(G107), .ZN(new_n230));
  OAI21_X1  g044(.A(G101), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT3), .B1(new_n229), .B2(G107), .ZN(new_n232));
  AOI21_X1  g046(.A(G101), .B1(new_n229), .B2(G107), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n227), .A3(G104), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n231), .A2(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n220), .A2(new_n226), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT78), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n220), .A2(KEYINPUT78), .A3(new_n237), .A4(new_n226), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n223), .B1(new_n243), .B2(KEYINPUT1), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n209), .A2(new_n210), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n221), .B1(new_n245), .B2(G146), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n226), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n237), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AND3_X1   g063(.A1(new_n242), .A2(KEYINPUT79), .A3(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT77), .ZN(new_n251));
  OR3_X1    g065(.A1(new_n251), .A2(KEYINPUT79), .A3(KEYINPUT12), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(new_n242), .B2(new_n249), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n206), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n242), .A2(new_n249), .ZN(new_n255));
  INV_X1    g069(.A(new_n206), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(new_n251), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(KEYINPUT12), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n254), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT10), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n247), .A2(new_n261), .A3(new_n248), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n237), .B1(new_n220), .B2(new_n226), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n262), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  NOR2_X1   g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n211), .B(new_n267), .C1(new_n218), .C2(new_n219), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n265), .B(new_n222), .C1(new_n225), .C2(new_n208), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n229), .A2(G107), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n232), .A2(new_n235), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT4), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G101), .ZN(new_n273));
  AND3_X1   g087(.A1(new_n268), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n236), .A2(KEYINPUT4), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT75), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n271), .A2(G101), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n276), .B1(new_n275), .B2(new_n277), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n274), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n264), .A2(new_n256), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(KEYINPUT76), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT76), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n264), .A2(new_n280), .A3(new_n283), .A4(new_n256), .ZN(new_n284));
  AND2_X1   g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n193), .B1(new_n260), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n193), .B1(new_n282), .B2(new_n284), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n264), .A2(new_n280), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n206), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G469), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n187), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n282), .A2(new_n284), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(new_n289), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n193), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n242), .A2(KEYINPUT79), .A3(new_n249), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n240), .A2(new_n241), .B1(new_n248), .B2(new_n247), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n297), .B1(new_n298), .B2(new_n252), .ZN(new_n299));
  AOI22_X1  g113(.A1(new_n299), .A2(new_n206), .B1(KEYINPUT12), .B2(new_n258), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT81), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n300), .B1(new_n287), .B2(new_n301), .ZN(new_n302));
  AOI211_X1 g116(.A(KEYINPUT81), .B(new_n193), .C1(new_n282), .C2(new_n284), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n296), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G902), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n292), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n192), .B1(new_n300), .B2(new_n294), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n294), .A2(new_n192), .A3(new_n289), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT80), .A3(G469), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n293), .A2(new_n306), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT9), .B(G234), .ZN(new_n312));
  OAI21_X1  g126(.A(G221), .B1(new_n312), .B2(G902), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G217), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(G234), .B2(new_n305), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n223), .B(G119), .C1(KEYINPUT71), .C2(KEYINPUT23), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT23), .ZN(new_n319));
  INV_X1    g133(.A(G119), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n319), .B1(new_n320), .B2(G128), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT71), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n320), .B2(G128), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n318), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G110), .ZN(new_n325));
  XOR2_X1   g139(.A(KEYINPUT24), .B(G110), .Z(new_n326));
  XNOR2_X1  g140(.A(G119), .B(G128), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g142(.A(G125), .B(G140), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT16), .ZN(new_n330));
  INV_X1    g144(.A(G140), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G125), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n332), .A2(KEYINPUT16), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n330), .A2(G146), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(G146), .B1(new_n330), .B2(new_n333), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n325), .B(new_n328), .C1(new_n335), .C2(new_n336), .ZN(new_n337));
  OAI22_X1  g151(.A1(new_n324), .A2(G110), .B1(new_n327), .B2(new_n326), .ZN(new_n338));
  INV_X1    g152(.A(G125), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G140), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n332), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n338), .B(new_n334), .C1(G146), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n344));
  XNOR2_X1  g158(.A(new_n344), .B(KEYINPUT72), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G137), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n337), .A2(new_n342), .A3(new_n347), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n349), .A2(new_n305), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n349), .A2(KEYINPUT25), .A3(new_n305), .A4(new_n350), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n317), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n349), .A2(new_n350), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n316), .A2(G902), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n357), .B(KEYINPUT73), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n320), .A2(G116), .ZN(new_n362));
  INV_X1    g176(.A(G116), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G119), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT68), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n362), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n365), .B1(new_n362), .B2(new_n364), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NOR2_X1   g182(.A1(KEYINPUT2), .A2(G113), .ZN(new_n369));
  NAND2_X1  g183(.A1(KEYINPUT2), .A2(G113), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(KEYINPUT67), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT67), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(KEYINPUT2), .A3(G113), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n369), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n368), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n371), .A2(new_n373), .ZN(new_n377));
  INV_X1    g191(.A(new_n369), .ZN(new_n378));
  XNOR2_X1  g192(.A(G116), .B(G119), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n377), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n376), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n220), .A2(new_n226), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n200), .A2(new_n201), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n197), .A2(G134), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(new_n199), .A3(G131), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT30), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n206), .A2(new_n268), .A3(new_n269), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n389), .B1(new_n388), .B2(new_n390), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n382), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(G237), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n188), .A3(G210), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n395), .B(KEYINPUT27), .ZN(new_n396));
  XNOR2_X1  g210(.A(KEYINPUT26), .B(G101), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n396), .B(new_n397), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n366), .A2(new_n374), .A3(new_n367), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(new_n380), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n388), .A2(new_n400), .A3(new_n390), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n393), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(KEYINPUT31), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT31), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n393), .A2(new_n404), .A3(new_n398), .A4(new_n401), .ZN(new_n405));
  AND3_X1   g219(.A1(new_n388), .A2(new_n400), .A3(new_n390), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n400), .B1(new_n388), .B2(new_n390), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT28), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT28), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n401), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n398), .B(KEYINPUT69), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n403), .A2(new_n405), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(G472), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n415), .A2(new_n416), .A3(new_n305), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT32), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT32), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n415), .A2(new_n419), .A3(new_n416), .A4(new_n305), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT70), .ZN(new_n422));
  NAND2_X1  g236(.A1(G472), .A2(G902), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT29), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n408), .A2(new_n424), .A3(new_n410), .A4(new_n412), .ZN(new_n425));
  INV_X1    g239(.A(new_n398), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n206), .A2(new_n268), .A3(new_n269), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n220), .A2(new_n226), .B1(new_n384), .B2(new_n386), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT30), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n388), .A2(new_n389), .A3(new_n390), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n400), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n426), .B1(new_n431), .B2(new_n406), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n425), .A2(new_n432), .A3(G472), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n382), .B1(new_n427), .B2(new_n428), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n409), .B1(new_n434), .B2(new_n401), .ZN(new_n435));
  INV_X1    g249(.A(new_n410), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n424), .B1(new_n437), .B2(new_n398), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n422), .B(new_n423), .C1(new_n433), .C2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n408), .A2(new_n398), .A3(new_n410), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT29), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n442), .A2(G472), .A3(new_n425), .A4(new_n432), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n422), .B1(new_n443), .B2(new_n423), .ZN(new_n444));
  NOR2_X1   g258(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n361), .B1(new_n421), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  XNOR2_X1  g261(.A(G110), .B(G122), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT5), .B1(new_n366), .B2(new_n367), .ZN(new_n450));
  OR2_X1    g264(.A1(new_n362), .A2(KEYINPUT5), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n451), .A2(G113), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n380), .B1(new_n450), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n277), .A2(KEYINPUT4), .A3(new_n236), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT75), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n273), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n376), .B2(new_n381), .ZN(new_n459));
  AOI221_X4 g273(.A(new_n449), .B1(new_n248), .B2(new_n453), .C1(new_n457), .C2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n339), .B1(new_n268), .B2(new_n269), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n220), .A2(new_n339), .A3(new_n226), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT82), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT82), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n220), .A2(new_n464), .A3(new_n339), .A4(new_n226), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n461), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(KEYINPUT85), .B(KEYINPUT7), .ZN(new_n467));
  XOR2_X1   g281(.A(KEYINPUT83), .B(G224), .Z(new_n468));
  AOI21_X1  g282(.A(new_n467), .B1(new_n468), .B2(new_n188), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n463), .A2(new_n465), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n468), .A2(new_n188), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(KEYINPUT7), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n461), .A2(new_n473), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NOR3_X1   g289(.A1(new_n460), .A2(new_n470), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n379), .A2(KEYINPUT5), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n452), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n478), .A2(new_n381), .A3(new_n248), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n453), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(new_n237), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT84), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n481), .A2(KEYINPUT84), .A3(new_n237), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n448), .B(KEYINPUT8), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n476), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n273), .B1(new_n399), .B2(new_n380), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n456), .B2(new_n455), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n453), .A2(new_n248), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n449), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n457), .A2(new_n459), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n492), .A3(new_n448), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(KEYINPUT6), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT6), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n498), .B(new_n449), .C1(new_n491), .C2(new_n493), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n466), .B(new_n472), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(G210), .B1(G237), .B2(G902), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n489), .A2(new_n501), .A3(new_n305), .A4(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(G902), .B1(new_n476), .B2(new_n488), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n502), .B1(new_n505), .B2(new_n501), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n447), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(G475), .A2(G902), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n394), .A2(new_n188), .A3(G214), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n216), .A3(new_n217), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n394), .A2(new_n188), .A3(G143), .A4(G214), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G131), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(KEYINPUT87), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n201), .A3(new_n511), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT17), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT87), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n512), .A2(new_n517), .A3(G131), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n514), .A2(new_n515), .A3(new_n516), .A4(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n335), .A2(new_n336), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n517), .B1(new_n512), .B2(G131), .ZN(new_n521));
  AOI211_X1 g335(.A(KEYINPUT87), .B(new_n201), .C1(new_n510), .C2(new_n511), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT17), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n519), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(G113), .B(G122), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT89), .B(G104), .ZN(new_n526));
  XOR2_X1   g340(.A(new_n525), .B(new_n526), .Z(new_n527));
  NAND2_X1  g341(.A1(KEYINPUT18), .A2(G131), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n510), .A2(new_n528), .A3(new_n511), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n512), .A2(KEYINPUT18), .A3(G131), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n329), .B(G146), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT86), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n329), .B(new_n208), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n534), .A2(KEYINPUT86), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n529), .B(new_n530), .C1(new_n533), .C2(new_n535), .ZN(new_n536));
  AND3_X1   g350(.A1(new_n524), .A2(new_n527), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n514), .A2(new_n518), .A3(new_n515), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT88), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n329), .A2(KEYINPUT19), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n332), .A2(new_n340), .A3(KEYINPUT19), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n539), .B1(new_n542), .B2(G146), .ZN(new_n543));
  OAI211_X1 g357(.A(KEYINPUT88), .B(new_n208), .C1(new_n540), .C2(new_n541), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n538), .A2(new_n334), .A3(new_n543), .A4(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n527), .B1(new_n545), .B2(new_n536), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n508), .B1(new_n537), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT20), .ZN(new_n548));
  INV_X1    g362(.A(new_n538), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n543), .A2(new_n334), .A3(new_n544), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n536), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n527), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n524), .A2(new_n527), .A3(new_n536), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT20), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n555), .A2(new_n556), .A3(new_n508), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n527), .B1(new_n524), .B2(new_n536), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n305), .B1(new_n537), .B2(new_n558), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n548), .A2(new_n557), .B1(G475), .B2(new_n559), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n312), .A2(new_n315), .A3(G953), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NOR3_X1   g376(.A1(new_n209), .A2(new_n210), .A3(new_n223), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n212), .A2(G128), .ZN(new_n564));
  OAI21_X1  g378(.A(KEYINPUT92), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n216), .A2(G128), .A3(new_n217), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT92), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n223), .A2(G143), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n565), .A2(new_n569), .A3(new_n195), .ZN(new_n570));
  XNOR2_X1  g384(.A(G116), .B(G122), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(new_n227), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n216), .A2(KEYINPUT13), .A3(G128), .A4(new_n217), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT13), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n564), .A2(new_n575), .ZN(new_n576));
  OAI211_X1 g390(.A(KEYINPUT90), .B(new_n574), .C1(new_n563), .C2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT90), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n566), .B(new_n578), .C1(new_n575), .C2(new_n564), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n577), .A2(G134), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT91), .ZN(new_n581));
  AOI22_X1  g395(.A1(new_n245), .A2(G128), .B1(KEYINPUT13), .B2(new_n568), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n195), .B1(new_n582), .B2(new_n578), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT91), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n577), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n573), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  OR2_X1    g400(.A1(new_n363), .A2(G122), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n227), .B1(new_n587), .B2(KEYINPUT14), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n588), .B(new_n571), .Z(new_n589));
  AOI21_X1  g403(.A(new_n195), .B1(new_n565), .B2(new_n569), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n591), .B2(new_n570), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n562), .B1(new_n586), .B2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n573), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n580), .A2(KEYINPUT91), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n584), .B1(new_n583), .B2(new_n577), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n588), .B(new_n571), .ZN(new_n598));
  INV_X1    g412(.A(new_n570), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n598), .B1(new_n599), .B2(new_n590), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n597), .A2(new_n600), .A3(new_n561), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n593), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(G478), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT93), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n604), .A2(KEYINPUT15), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(KEYINPUT15), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n603), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n602), .B(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(G952), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n610), .A2(KEYINPUT94), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n610), .A2(KEYINPUT94), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n188), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n613), .B1(G234), .B2(G237), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT21), .B(G898), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n305), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n560), .A2(new_n609), .A3(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n507), .A2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n314), .A2(new_n446), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT95), .B(G101), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G3));
  OAI211_X1 g437(.A(new_n447), .B(new_n618), .C1(new_n504), .C2(new_n506), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n586), .A2(new_n592), .A3(new_n562), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n561), .B1(new_n597), .B2(new_n600), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT33), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT33), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n593), .A2(new_n601), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n627), .A2(G478), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n603), .A2(new_n305), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n602), .B2(new_n603), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n560), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n624), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n415), .A2(new_n305), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(G472), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n417), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n361), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n314), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT34), .B(G104), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G6));
  NAND2_X1  g457(.A1(new_n559), .A2(G475), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n556), .B1(new_n555), .B2(new_n508), .ZN(new_n645));
  INV_X1    g459(.A(new_n508), .ZN(new_n646));
  AOI211_X1 g460(.A(KEYINPUT20), .B(new_n646), .C1(new_n553), .C2(new_n554), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n644), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n648), .A2(new_n609), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n624), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n314), .A2(new_n640), .A3(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  INV_X1    g467(.A(new_n355), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n348), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(new_n343), .ZN(new_n656));
  INV_X1    g470(.A(new_n358), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n638), .A2(new_n417), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(KEYINPUT96), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n314), .A2(new_n620), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT37), .B(G110), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G12));
  OAI211_X1 g478(.A(new_n447), .B(new_n659), .C1(new_n504), .C2(new_n506), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n421), .B2(new_n445), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n614), .B1(new_n667), .B2(new_n616), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n649), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n666), .A2(new_n311), .A3(new_n313), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  INV_X1    g485(.A(new_n402), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n412), .B1(new_n401), .B2(new_n434), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n305), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(G472), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n421), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(new_n676), .B(KEYINPUT97), .Z(new_n677));
  NOR2_X1   g491(.A1(new_n560), .A2(new_n609), .ZN(new_n678));
  INV_X1    g492(.A(new_n659), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n678), .A2(new_n447), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT98), .ZN(new_n681));
  AND2_X1   g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n502), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n497), .A2(new_n499), .A3(new_n500), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n471), .A2(new_n474), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n496), .B(new_n685), .C1(new_n466), .C2(new_n469), .ZN(new_n686));
  INV_X1    g500(.A(new_n487), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n484), .B2(new_n485), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n305), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n683), .B1(new_n684), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n503), .ZN(new_n691));
  XOR2_X1   g505(.A(new_n691), .B(KEYINPUT38), .Z(new_n692));
  NOR2_X1   g506(.A1(new_n680), .A2(new_n681), .ZN(new_n693));
  NOR4_X1   g507(.A1(new_n677), .A2(new_n682), .A3(new_n692), .A4(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(new_n668), .B(KEYINPUT39), .Z(new_n695));
  NAND2_X1  g509(.A1(new_n314), .A2(new_n695), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(KEYINPUT40), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n694), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(new_n225), .ZN(G45));
  INV_X1    g514(.A(new_n668), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n634), .A2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n666), .A2(new_n311), .A3(new_n313), .A4(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G146), .ZN(G48));
  AND3_X1   g519(.A1(new_n304), .A2(new_n292), .A3(new_n305), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n292), .B1(new_n304), .B2(new_n305), .ZN(new_n707));
  INV_X1    g521(.A(new_n313), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n706), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n446), .A3(new_n636), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT41), .B(G113), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G15));
  NAND3_X1  g526(.A1(new_n709), .A2(new_n446), .A3(new_n650), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G116), .ZN(G18));
  NAND4_X1  g528(.A1(new_n560), .A2(new_n659), .A3(new_n609), .A4(new_n618), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n421), .B2(new_n445), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n706), .A2(new_n707), .ZN(new_n717));
  INV_X1    g531(.A(new_n447), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n690), .B2(new_n503), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n716), .A2(new_n717), .A3(new_n313), .A4(new_n719), .ZN(new_n720));
  XOR2_X1   g534(.A(KEYINPUT99), .B(G119), .Z(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G21));
  NAND3_X1  g536(.A1(new_n719), .A2(new_n678), .A3(new_n618), .ZN(new_n723));
  OR3_X1    g537(.A1(new_n355), .A2(KEYINPUT100), .A3(new_n359), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT100), .B1(new_n355), .B2(new_n359), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n638), .A3(new_n417), .ZN(new_n727));
  NOR2_X1   g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n709), .ZN(new_n729));
  XNOR2_X1  g543(.A(KEYINPUT101), .B(G122), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G24));
  NOR2_X1   g545(.A1(new_n702), .A2(new_n660), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n709), .A2(new_n719), .A3(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G125), .ZN(G27));
  INV_X1    g548(.A(KEYINPUT42), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT103), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n690), .A2(new_n447), .A3(new_n503), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT102), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT102), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n690), .A2(new_n739), .A3(new_n447), .A4(new_n503), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n738), .A2(new_n313), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n309), .A2(G469), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n306), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n736), .B1(new_n741), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n738), .A2(new_n313), .A3(new_n740), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n306), .A2(new_n742), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n745), .A2(new_n746), .A3(KEYINPUT103), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n446), .B(new_n703), .C1(new_n744), .C2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT104), .ZN(new_n749));
  AOI22_X1  g563(.A1(new_n402), .A2(KEYINPUT31), .B1(new_n411), .B2(new_n413), .ZN(new_n750));
  AOI21_X1  g564(.A(G902), .B1(new_n750), .B2(new_n405), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n419), .B1(new_n751), .B2(new_n416), .ZN(new_n752));
  INV_X1    g566(.A(new_n420), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n749), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n418), .A2(KEYINPUT104), .A3(new_n420), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n445), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n726), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT105), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(KEYINPUT105), .A3(new_n726), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n703), .A2(KEYINPUT42), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n741), .A2(new_n736), .A3(new_n743), .ZN(new_n763));
  OAI21_X1  g577(.A(KEYINPUT103), .B1(new_n745), .B2(new_n746), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n735), .A2(new_n748), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(new_n201), .ZN(G33));
  OAI211_X1 g581(.A(new_n446), .B(new_n669), .C1(new_n744), .C2(new_n747), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G134), .ZN(G36));
  NAND2_X1  g583(.A1(new_n738), .A2(new_n740), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(KEYINPUT106), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n648), .A2(new_n633), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT43), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n773), .A2(new_n639), .A3(new_n659), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n771), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n774), .A2(new_n775), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT107), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n781));
  OAI21_X1  g595(.A(new_n781), .B1(new_n307), .B2(new_n308), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n286), .A2(KEYINPUT45), .A3(new_n290), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n783), .A3(G469), .ZN(new_n784));
  NAND2_X1  g598(.A1(G469), .A2(G902), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT46), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n706), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n785), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n708), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n789), .A2(new_n695), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n776), .A2(KEYINPUT107), .A3(new_n777), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n780), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G137), .ZN(G39));
  NOR2_X1   g607(.A1(KEYINPUT108), .A2(KEYINPUT47), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n789), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n795), .B1(new_n789), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n421), .A2(new_n445), .ZN(new_n798));
  NOR4_X1   g612(.A1(new_n770), .A2(new_n798), .A3(new_n360), .A4(new_n702), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G140), .ZN(G42));
  NOR2_X1   g615(.A1(new_n708), .A2(new_n718), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n692), .A2(new_n726), .A3(new_n772), .A4(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n717), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n803), .B1(KEYINPUT49), .B2(new_n804), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n805), .B(new_n677), .C1(KEYINPUT49), .C2(new_n804), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n741), .A2(new_n614), .A3(new_n717), .ZN(new_n807));
  AND3_X1   g621(.A1(new_n677), .A2(new_n360), .A3(new_n807), .ZN(new_n808));
  XOR2_X1   g622(.A(new_n808), .B(KEYINPUT116), .Z(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n634), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n761), .A2(new_n773), .A3(new_n807), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT48), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n812), .A2(KEYINPUT118), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n812), .A2(KEYINPUT118), .ZN(new_n814));
  OR3_X1    g628(.A1(new_n811), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n727), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n773), .A2(new_n614), .A3(new_n816), .ZN(new_n817));
  NOR4_X1   g631(.A1(new_n817), .A2(new_n804), .A3(new_n708), .A4(new_n507), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n818), .A2(new_n613), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n811), .A2(new_n813), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n810), .A2(new_n815), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n692), .A2(new_n718), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n817), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n823), .A2(KEYINPUT50), .A3(new_n709), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT50), .B1(new_n823), .B2(new_n709), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n807), .A2(new_n773), .ZN(new_n826));
  OAI22_X1  g640(.A1(new_n824), .A2(new_n825), .B1(new_n660), .B2(new_n826), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n560), .A2(new_n633), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n809), .A2(KEYINPUT117), .A3(new_n828), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n808), .A2(KEYINPUT116), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n808), .A2(KEYINPUT116), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n827), .B1(new_n829), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n771), .A2(new_n817), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n804), .A2(new_n313), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n836), .B1(new_n797), .B2(new_n837), .ZN(new_n838));
  AND2_X1   g652(.A1(new_n838), .A2(KEYINPUT51), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n821), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  OR2_X1    g654(.A1(new_n797), .A2(KEYINPUT115), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n797), .A2(KEYINPUT115), .ZN(new_n842));
  OAI211_X1 g656(.A(new_n841), .B(new_n842), .C1(new_n313), .C2(new_n804), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n836), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n835), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n840), .B1(new_n845), .B2(KEYINPUT51), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT112), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n560), .A2(new_n609), .A3(new_n848), .A4(new_n701), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n305), .B1(new_n625), .B2(new_n626), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n608), .ZN(new_n851));
  INV_X1    g665(.A(new_n608), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n602), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n853), .A3(new_n701), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT112), .B1(new_n648), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n679), .B1(new_n849), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n798), .A2(new_n856), .A3(new_n740), .A4(new_n738), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n311), .A2(new_n313), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n763), .A2(new_n764), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n859), .B1(new_n860), .B2(new_n732), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n710), .A2(new_n713), .A3(new_n720), .A4(new_n729), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n861), .A2(new_n768), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT111), .ZN(new_n864));
  OAI21_X1  g678(.A(KEYINPUT110), .B1(new_n624), .B2(new_n649), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT109), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n866), .B1(new_n560), .B2(new_n633), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n648), .A2(KEYINPUT109), .A3(new_n630), .A4(new_n632), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n867), .A2(new_n868), .A3(new_n719), .A4(new_n618), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n648), .A2(new_n609), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT110), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n719), .A2(new_n870), .A3(new_n871), .A4(new_n618), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n865), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n311), .A2(new_n313), .A3(new_n640), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n311), .A2(new_n313), .A3(new_n620), .ZN(new_n877));
  INV_X1    g691(.A(new_n446), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT96), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n660), .B(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n877), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n864), .B1(new_n876), .B2(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n314), .A2(new_n640), .A3(new_n873), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n621), .A2(new_n662), .A3(new_n883), .A4(KEYINPUT111), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n748), .A2(new_n735), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n761), .A2(new_n765), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n314), .B(new_n666), .C1(new_n669), .C2(new_n703), .ZN(new_n889));
  OR3_X1    g703(.A1(new_n659), .A2(KEYINPUT113), .A3(new_n668), .ZN(new_n890));
  OAI21_X1  g704(.A(KEYINPUT113), .B1(new_n659), .B2(new_n668), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n708), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n719), .A2(new_n678), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n676), .A3(new_n893), .A4(new_n743), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n889), .A2(KEYINPUT52), .A3(new_n733), .A4(new_n894), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n670), .A2(new_n704), .A3(new_n733), .A4(new_n894), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT52), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n863), .A2(new_n885), .A3(new_n888), .A4(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT53), .ZN(new_n901));
  OR2_X1    g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n732), .B1(new_n744), .B2(new_n747), .ZN(new_n903));
  INV_X1    g717(.A(new_n859), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n862), .A2(new_n768), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n766), .A2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT114), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n896), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(KEYINPUT52), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n896), .A2(new_n907), .A3(new_n897), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n906), .A2(new_n885), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n901), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n847), .B1(new_n902), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n900), .A2(new_n901), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n906), .A2(KEYINPUT53), .A3(new_n885), .A4(new_n911), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(KEYINPUT54), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n846), .A2(new_n914), .A3(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(G952), .A2(G953), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n806), .B1(new_n919), .B2(new_n920), .ZN(G75));
  NOR2_X1   g735(.A1(new_n188), .A2(G952), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n305), .B1(new_n915), .B2(new_n916), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT56), .B1(new_n924), .B2(G210), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n497), .A2(new_n499), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(new_n500), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT55), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n923), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT56), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n917), .A2(G902), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT119), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n924), .A2(KEYINPUT119), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n936), .A2(new_n502), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT120), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n931), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT120), .B1(new_n936), .B2(new_n502), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n929), .B1(new_n939), .B2(new_n940), .ZN(G51));
  OR2_X1    g755(.A1(new_n936), .A2(new_n784), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n917), .B(new_n847), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n785), .B(KEYINPUT57), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n304), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n922), .B1(new_n942), .B2(new_n945), .ZN(G54));
  AND2_X1   g760(.A1(KEYINPUT58), .A2(G475), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n934), .A2(new_n935), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n555), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n948), .A2(KEYINPUT122), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT119), .B1(new_n917), .B2(G902), .ZN(new_n951));
  AOI211_X1 g765(.A(new_n933), .B(new_n305), .C1(new_n915), .C2(new_n916), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n555), .A2(new_n947), .ZN(new_n954));
  AOI21_X1  g768(.A(KEYINPUT121), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AND4_X1   g769(.A1(KEYINPUT121), .A2(new_n934), .A3(new_n935), .A4(new_n954), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n950), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n555), .B1(new_n953), .B2(new_n947), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n923), .B1(new_n958), .B2(KEYINPUT122), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n957), .A2(new_n959), .ZN(G60));
  AND2_X1   g774(.A1(new_n627), .A2(new_n629), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n631), .B(KEYINPUT59), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n923), .B1(new_n943), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT123), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n967), .B(new_n923), .C1(new_n943), .C2(new_n964), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n914), .A2(new_n918), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n961), .B1(new_n969), .B2(new_n962), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n966), .A2(new_n968), .A3(new_n970), .ZN(G63));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n972));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT60), .Z(new_n974));
  AND2_X1   g788(.A1(new_n917), .A2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n922), .B1(new_n975), .B2(new_n656), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n917), .A2(new_n974), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(new_n356), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n972), .B1(new_n976), .B2(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(G66));
  INV_X1    g795(.A(new_n615), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n188), .B1(new_n982), .B2(new_n468), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n885), .A2(new_n862), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n983), .B1(new_n984), .B2(new_n188), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n926), .B1(G898), .B2(new_n188), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n985), .B(new_n986), .Z(G69));
  AOI21_X1  g801(.A(new_n870), .B1(new_n867), .B2(new_n868), .ZN(new_n988));
  OR4_X1    g802(.A1(new_n878), .A2(new_n696), .A3(new_n770), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n792), .A2(new_n989), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT125), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n889), .A2(new_n733), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n699), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(KEYINPUT62), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n800), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n188), .B1(new_n992), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n429), .A2(new_n430), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(new_n542), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1000), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n993), .A2(new_n768), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n792), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n790), .A2(new_n761), .A3(new_n893), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n800), .A2(new_n1005), .ZN(new_n1006));
  NAND4_X1  g820(.A1(new_n1004), .A2(KEYINPUT127), .A3(new_n1006), .A4(new_n888), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT127), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n792), .A2(new_n800), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1008), .B1(new_n1009), .B2(new_n766), .ZN(new_n1010));
  AOI21_X1  g824(.A(G953), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n188), .A2(G900), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT126), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1002), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1015));
  AND3_X1   g829(.A1(new_n1001), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1015), .B1(new_n1001), .B2(new_n1014), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1016), .A2(new_n1017), .ZN(G72));
  NOR2_X1   g832(.A1(new_n431), .A2(new_n406), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n984), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1007), .A2(new_n1010), .A3(new_n1021), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n423), .B(KEYINPUT63), .Z(new_n1023));
  AOI211_X1 g837(.A(new_n398), .B(new_n1020), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1020), .A2(new_n398), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n990), .B(KEYINPUT125), .ZN(new_n1026));
  NAND4_X1  g840(.A1(new_n1026), .A2(new_n800), .A3(new_n1021), .A4(new_n996), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1025), .B1(new_n1027), .B2(new_n1023), .ZN(new_n1028));
  INV_X1    g842(.A(new_n432), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1023), .B1(new_n1029), .B2(new_n672), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1030), .B1(new_n902), .B2(new_n913), .ZN(new_n1031));
  NOR4_X1   g845(.A1(new_n1024), .A2(new_n1028), .A3(new_n922), .A4(new_n1031), .ZN(G57));
endmodule


