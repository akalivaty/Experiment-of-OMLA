

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731;

  AND2_X1 U366 ( .A1(n613), .A2(n612), .ZN(n672) );
  XNOR2_X1 U367 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U368 ( .A(n465), .B(n390), .ZN(n716) );
  AND2_X1 U369 ( .A1(n366), .A2(n367), .ZN(n640) );
  XNOR2_X2 U370 ( .A(n595), .B(KEYINPUT1), .ZN(n578) );
  XNOR2_X2 U371 ( .A(n499), .B(KEYINPUT0), .ZN(n571) );
  NOR2_X1 U372 ( .A1(n703), .A2(n718), .ZN(n642) );
  NOR2_X1 U373 ( .A1(n634), .A2(n633), .ZN(n635) );
  OR2_X1 U374 ( .A1(n642), .A2(n344), .ZN(n356) );
  XNOR2_X1 U375 ( .A(n371), .B(n352), .ZN(n703) );
  AND2_X1 U376 ( .A1(n370), .A2(KEYINPUT44), .ZN(n353) );
  XNOR2_X1 U377 ( .A(n562), .B(KEYINPUT67), .ZN(n366) );
  XNOR2_X1 U378 ( .A(n373), .B(n351), .ZN(n639) );
  NAND2_X1 U379 ( .A1(n375), .A2(n374), .ZN(n373) );
  INV_X1 U380 ( .A(n564), .ZN(n374) );
  NAND2_X1 U381 ( .A1(n384), .A2(n381), .ZN(n613) );
  AND2_X1 U382 ( .A1(n386), .A2(n347), .ZN(n384) );
  XNOR2_X1 U383 ( .A(n458), .B(n457), .ZN(n688) );
  XNOR2_X1 U384 ( .A(n452), .B(n451), .ZN(n458) );
  XNOR2_X1 U385 ( .A(n411), .B(n410), .ZN(n461) );
  XNOR2_X1 U386 ( .A(n456), .B(n350), .ZN(n457) );
  NOR2_X1 U387 ( .A1(n624), .A2(n589), .ZN(n590) );
  NOR2_X2 U388 ( .A1(n570), .A2(n445), .ZN(n586) );
  XNOR2_X2 U389 ( .A(n589), .B(n507), .ZN(n663) );
  NOR2_X1 U390 ( .A1(n581), .A2(KEYINPUT44), .ZN(n365) );
  NAND2_X1 U391 ( .A1(n566), .A2(n567), .ZN(n368) );
  NAND2_X1 U392 ( .A1(n719), .A2(G234), .ZN(n411) );
  AND2_X1 U393 ( .A1(n630), .A2(KEYINPUT2), .ZN(n357) );
  INV_X1 U394 ( .A(KEYINPUT19), .ZN(n385) );
  INV_X1 U395 ( .A(n493), .ZN(n383) );
  XNOR2_X1 U396 ( .A(n428), .B(n427), .ZN(n648) );
  NAND2_X1 U397 ( .A1(n361), .A2(n644), .ZN(n359) );
  XNOR2_X1 U398 ( .A(n588), .B(n587), .ZN(n624) );
  BUF_X1 U399 ( .A(n523), .Z(n517) );
  AND2_X1 U400 ( .A1(n380), .A2(n379), .ZN(n577) );
  INV_X1 U401 ( .A(n519), .ZN(n379) );
  OR2_X1 U402 ( .A1(n719), .A2(G952), .ZN(n659) );
  XNOR2_X1 U403 ( .A(n511), .B(KEYINPUT72), .ZN(n591) );
  AND2_X1 U404 ( .A1(n510), .A2(n529), .ZN(n511) );
  NAND2_X1 U405 ( .A1(n366), .A2(n365), .ZN(n364) );
  AND2_X1 U406 ( .A1(n583), .A2(n662), .ZN(n355) );
  NOR2_X1 U407 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U408 ( .A(n470), .B(n404), .ZN(n405) );
  XNOR2_X1 U409 ( .A(KEYINPUT10), .B(KEYINPUT71), .ZN(n404) );
  NOR2_X1 U410 ( .A1(n505), .A2(n500), .ZN(n389) );
  AND2_X1 U411 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U412 ( .A(G119), .B(G113), .ZN(n425) );
  XNOR2_X1 U413 ( .A(KEYINPUT73), .B(KEYINPUT3), .ZN(n424) );
  XNOR2_X1 U414 ( .A(G119), .B(G128), .ZN(n407) );
  XOR2_X1 U415 ( .A(KEYINPUT101), .B(G107), .Z(n464) );
  XOR2_X1 U416 ( .A(G140), .B(G104), .Z(n454) );
  XNOR2_X1 U417 ( .A(n716), .B(n392), .ZN(n428) );
  XNOR2_X1 U418 ( .A(G107), .B(G104), .ZN(n394) );
  XNOR2_X1 U419 ( .A(KEYINPUT77), .B(G110), .ZN(n393) );
  INV_X1 U420 ( .A(KEYINPUT78), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n522), .B(n521), .ZN(n563) );
  INV_X1 U422 ( .A(KEYINPUT33), .ZN(n521) );
  NOR2_X1 U423 ( .A1(n520), .A2(n578), .ZN(n522) );
  XNOR2_X1 U424 ( .A(n377), .B(n376), .ZN(n375) );
  INV_X1 U425 ( .A(KEYINPUT34), .ZN(n376) );
  NAND2_X1 U426 ( .A1(n563), .A2(n568), .ZN(n377) );
  NOR2_X1 U427 ( .A1(n542), .A2(KEYINPUT19), .ZN(n382) );
  OR2_X1 U428 ( .A1(n595), .A2(n525), .ZN(n570) );
  INV_X1 U429 ( .A(KEYINPUT64), .ZN(n395) );
  INV_X1 U430 ( .A(G953), .ZN(n636) );
  INV_X1 U431 ( .A(KEYINPUT109), .ZN(n515) );
  NAND2_X1 U432 ( .A1(n577), .A2(n503), .ZN(n378) );
  XNOR2_X1 U433 ( .A(n569), .B(KEYINPUT31), .ZN(n678) );
  OR2_X1 U434 ( .A1(n646), .A2(n641), .ZN(n344) );
  NOR2_X1 U435 ( .A1(n572), .A2(n571), .ZN(n345) );
  AND2_X1 U436 ( .A1(n383), .A2(n387), .ZN(n346) );
  OR2_X1 U437 ( .A1(n387), .A2(n385), .ZN(n347) );
  NOR2_X1 U438 ( .A1(n578), .A2(n526), .ZN(n348) );
  AND2_X1 U439 ( .A1(n368), .A2(n364), .ZN(n349) );
  INV_X1 U440 ( .A(n581), .ZN(n367) );
  AND2_X1 U441 ( .A1(G214), .A2(n455), .ZN(n350) );
  INV_X1 U442 ( .A(n542), .ZN(n387) );
  XOR2_X1 U443 ( .A(KEYINPUT80), .B(KEYINPUT35), .Z(n351) );
  XOR2_X1 U444 ( .A(n584), .B(KEYINPUT65), .Z(n352) );
  NAND2_X1 U445 ( .A1(n354), .A2(n353), .ZN(n369) );
  INV_X1 U446 ( .A(n640), .ZN(n354) );
  NOR2_X1 U447 ( .A1(n698), .A2(G902), .ZN(n419) );
  XNOR2_X1 U448 ( .A(n415), .B(n414), .ZN(n698) );
  NAND2_X1 U449 ( .A1(n372), .A2(n355), .ZN(n371) );
  NAND2_X2 U450 ( .A1(n356), .A2(n359), .ZN(n360) );
  NAND2_X1 U451 ( .A1(n358), .A2(n357), .ZN(n363) );
  INV_X1 U452 ( .A(n703), .ZN(n358) );
  NOR2_X4 U453 ( .A1(n647), .A2(n360), .ZN(n693) );
  INV_X1 U454 ( .A(n646), .ZN(n361) );
  XNOR2_X2 U455 ( .A(n363), .B(n362), .ZN(n647) );
  NAND2_X1 U456 ( .A1(n383), .A2(n382), .ZN(n381) );
  INV_X2 U457 ( .A(n405), .ZN(n450) );
  NAND2_X1 U458 ( .A1(n369), .A2(n349), .ZN(n372) );
  INV_X1 U459 ( .A(n566), .ZN(n370) );
  XNOR2_X2 U460 ( .A(n474), .B(G134), .ZN(n465) );
  XNOR2_X2 U461 ( .A(G143), .B(G128), .ZN(n474) );
  XNOR2_X2 U462 ( .A(n378), .B(n504), .ZN(n565) );
  XNOR2_X1 U463 ( .A(n557), .B(KEYINPUT22), .ZN(n380) );
  NAND2_X1 U464 ( .A1(n493), .A2(KEYINPUT19), .ZN(n386) );
  XNOR2_X2 U465 ( .A(n388), .B(n491), .ZN(n493) );
  NAND2_X1 U466 ( .A1(n680), .A2(n644), .ZN(n388) );
  NAND2_X1 U467 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U468 ( .A(n603), .B(KEYINPUT46), .ZN(n611) );
  XNOR2_X1 U469 ( .A(KEYINPUT4), .B(G131), .ZN(n390) );
  INV_X1 U470 ( .A(KEYINPUT8), .ZN(n410) );
  AND2_X1 U471 ( .A1(n604), .A2(n387), .ZN(n512) );
  BUF_X1 U472 ( .A(n598), .Z(n537) );
  INV_X1 U473 ( .A(KEYINPUT39), .ZN(n587) );
  BUF_X1 U474 ( .A(n693), .Z(n697) );
  XNOR2_X1 U475 ( .A(n524), .B(KEYINPUT41), .ZN(n598) );
  XNOR2_X1 U476 ( .A(n600), .B(n599), .ZN(n726) );
  XNOR2_X2 U477 ( .A(G101), .B(KEYINPUT70), .ZN(n391) );
  XNOR2_X2 U478 ( .A(n391), .B(KEYINPUT69), .ZN(n471) );
  XNOR2_X1 U479 ( .A(n471), .B(G146), .ZN(n392) );
  XOR2_X1 U480 ( .A(G137), .B(G140), .Z(n406) );
  XNOR2_X1 U481 ( .A(n394), .B(n393), .ZN(n482) );
  XNOR2_X2 U482 ( .A(n395), .B(G953), .ZN(n719) );
  AND2_X1 U483 ( .A1(n719), .A2(G227), .ZN(n396) );
  XNOR2_X1 U484 ( .A(n482), .B(n396), .ZN(n397) );
  XNOR2_X1 U485 ( .A(n406), .B(n397), .ZN(n398) );
  XNOR2_X1 U486 ( .A(n428), .B(n398), .ZN(n656) );
  INV_X1 U487 ( .A(G902), .ZN(n429) );
  NAND2_X1 U488 ( .A1(n656), .A2(n429), .ZN(n400) );
  INV_X1 U489 ( .A(G469), .ZN(n399) );
  XNOR2_X1 U490 ( .A(n400), .B(n399), .ZN(n595) );
  XOR2_X1 U491 ( .A(KEYINPUT20), .B(KEYINPUT95), .Z(n402) );
  XNOR2_X1 U492 ( .A(KEYINPUT15), .B(G902), .ZN(n644) );
  NAND2_X1 U493 ( .A1(G234), .A2(n644), .ZN(n401) );
  XNOR2_X1 U494 ( .A(n402), .B(n401), .ZN(n416) );
  NAND2_X1 U495 ( .A1(n416), .A2(G221), .ZN(n403) );
  XOR2_X1 U496 ( .A(KEYINPUT21), .B(n403), .Z(n529) );
  XOR2_X2 U497 ( .A(G146), .B(G125), .Z(n470) );
  XNOR2_X2 U498 ( .A(n406), .B(n450), .ZN(n715) );
  XOR2_X1 U499 ( .A(KEYINPUT94), .B(G110), .Z(n408) );
  XNOR2_X1 U500 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U501 ( .A(n715), .B(n409), .ZN(n415) );
  XOR2_X1 U502 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n413) );
  NAND2_X1 U503 ( .A1(G221), .A2(n461), .ZN(n412) );
  XNOR2_X1 U504 ( .A(n413), .B(n412), .ZN(n414) );
  NAND2_X1 U505 ( .A1(G217), .A2(n416), .ZN(n417) );
  XNOR2_X1 U506 ( .A(KEYINPUT25), .B(n417), .ZN(n418) );
  XNOR2_X1 U507 ( .A(n419), .B(n418), .ZN(n508) );
  NAND2_X1 U508 ( .A1(n529), .A2(n508), .ZN(n525) );
  XOR2_X1 U509 ( .A(KEYINPUT5), .B(KEYINPUT76), .Z(n421) );
  XNOR2_X1 U510 ( .A(G116), .B(G137), .ZN(n420) );
  XNOR2_X1 U511 ( .A(n421), .B(n420), .ZN(n423) );
  NOR2_X1 U512 ( .A1(G953), .A2(G237), .ZN(n455) );
  NAND2_X1 U513 ( .A1(n455), .A2(G210), .ZN(n422) );
  XNOR2_X1 U514 ( .A(n423), .B(n422), .ZN(n426) );
  XNOR2_X1 U515 ( .A(n425), .B(n424), .ZN(n481) );
  XNOR2_X1 U516 ( .A(n426), .B(n481), .ZN(n427) );
  NAND2_X1 U517 ( .A1(n648), .A2(n429), .ZN(n432) );
  INV_X1 U518 ( .A(KEYINPUT74), .ZN(n430) );
  XNOR2_X1 U519 ( .A(n430), .B(G472), .ZN(n431) );
  XNOR2_X2 U520 ( .A(n432), .B(n431), .ZN(n560) );
  OR2_X1 U521 ( .A1(G237), .A2(G902), .ZN(n488) );
  NAND2_X1 U522 ( .A1(G214), .A2(n488), .ZN(n433) );
  XNOR2_X1 U523 ( .A(n433), .B(KEYINPUT93), .ZN(n542) );
  NOR2_X1 U524 ( .A1(n560), .A2(n542), .ZN(n434) );
  XNOR2_X1 U525 ( .A(n434), .B(KEYINPUT30), .ZN(n444) );
  NAND2_X1 U526 ( .A1(G234), .A2(G237), .ZN(n436) );
  INV_X1 U527 ( .A(KEYINPUT14), .ZN(n435) );
  XNOR2_X1 U528 ( .A(n436), .B(n435), .ZN(n553) );
  INV_X1 U529 ( .A(n553), .ZN(n496) );
  NAND2_X1 U530 ( .A1(G902), .A2(n496), .ZN(n437) );
  NOR2_X1 U531 ( .A1(n719), .A2(n437), .ZN(n438) );
  XNOR2_X1 U532 ( .A(n438), .B(KEYINPUT107), .ZN(n439) );
  NOR2_X1 U533 ( .A1(G900), .A2(n439), .ZN(n440) );
  XNOR2_X1 U534 ( .A(n440), .B(KEYINPUT108), .ZN(n442) );
  NAND2_X1 U535 ( .A1(n636), .A2(G952), .ZN(n494) );
  NOR2_X1 U536 ( .A1(n553), .A2(n494), .ZN(n441) );
  NOR2_X1 U537 ( .A1(n442), .A2(n441), .ZN(n509) );
  INV_X1 U538 ( .A(n509), .ZN(n443) );
  NAND2_X1 U539 ( .A1(n444), .A2(n443), .ZN(n445) );
  XOR2_X1 U540 ( .A(KEYINPUT11), .B(KEYINPUT99), .Z(n447) );
  XNOR2_X1 U541 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n446) );
  XNOR2_X1 U542 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U543 ( .A(n448), .B(KEYINPUT12), .Z(n452) );
  XNOR2_X1 U544 ( .A(G143), .B(G122), .ZN(n449) );
  XNOR2_X1 U545 ( .A(G113), .B(G131), .ZN(n453) );
  XNOR2_X1 U546 ( .A(n454), .B(n453), .ZN(n456) );
  NOR2_X1 U547 ( .A1(G902), .A2(n688), .ZN(n460) );
  XNOR2_X1 U548 ( .A(KEYINPUT13), .B(G475), .ZN(n459) );
  XNOR2_X1 U549 ( .A(n460), .B(n459), .ZN(n505) );
  NAND2_X1 U550 ( .A1(G217), .A2(n461), .ZN(n463) );
  XOR2_X1 U551 ( .A(KEYINPUT9), .B(KEYINPUT7), .Z(n462) );
  XNOR2_X1 U552 ( .A(n463), .B(n462), .ZN(n468) );
  XNOR2_X1 U553 ( .A(G122), .B(G116), .ZN(n484) );
  XNOR2_X1 U554 ( .A(n464), .B(n484), .ZN(n466) );
  XOR2_X1 U555 ( .A(n466), .B(n465), .Z(n467) );
  XNOR2_X1 U556 ( .A(n468), .B(n467), .ZN(n694) );
  NOR2_X1 U557 ( .A1(G902), .A2(n694), .ZN(n469) );
  XNOR2_X1 U558 ( .A(n469), .B(G478), .ZN(n539) );
  INV_X1 U559 ( .A(n539), .ZN(n500) );
  NAND2_X1 U560 ( .A1(n505), .A2(n500), .ZN(n564) );
  XNOR2_X1 U561 ( .A(n471), .B(n470), .ZN(n476) );
  XNOR2_X1 U562 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n472) );
  XNOR2_X1 U563 ( .A(n472), .B(KEYINPUT90), .ZN(n473) );
  XNOR2_X1 U564 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U565 ( .A(n476), .B(n475), .ZN(n480) );
  XOR2_X1 U566 ( .A(KEYINPUT4), .B(KEYINPUT79), .Z(n478) );
  NAND2_X1 U567 ( .A1(G224), .A2(n719), .ZN(n477) );
  XNOR2_X1 U568 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U569 ( .A(n480), .B(n479), .ZN(n487) );
  XNOR2_X1 U570 ( .A(n482), .B(n481), .ZN(n486) );
  XNOR2_X1 U571 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n483) );
  XNOR2_X1 U572 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U573 ( .A(n486), .B(n485), .ZN(n710) );
  XNOR2_X1 U574 ( .A(n487), .B(n710), .ZN(n680) );
  XNOR2_X1 U575 ( .A(KEYINPUT91), .B(KEYINPUT92), .ZN(n490) );
  AND2_X1 U576 ( .A1(G210), .A2(n488), .ZN(n489) );
  XNOR2_X1 U577 ( .A(n490), .B(n489), .ZN(n491) );
  BUF_X1 U578 ( .A(n493), .Z(n523) );
  NOR2_X1 U579 ( .A1(n564), .A2(n517), .ZN(n492) );
  NAND2_X1 U580 ( .A1(n586), .A2(n492), .ZN(n616) );
  XNOR2_X1 U581 ( .A(n616), .B(G143), .ZN(G45) );
  NOR2_X1 U582 ( .A1(G898), .A2(n636), .ZN(n711) );
  NAND2_X1 U583 ( .A1(n711), .A2(G902), .ZN(n495) );
  NAND2_X1 U584 ( .A1(n495), .A2(n494), .ZN(n497) );
  AND2_X1 U585 ( .A1(n497), .A2(n496), .ZN(n498) );
  NAND2_X1 U586 ( .A1(n613), .A2(n498), .ZN(n499) );
  NAND2_X1 U587 ( .A1(n389), .A2(n529), .ZN(n501) );
  NOR2_X2 U588 ( .A1(n571), .A2(n501), .ZN(n557) );
  XNOR2_X1 U589 ( .A(n560), .B(KEYINPUT6), .ZN(n519) );
  BUF_X1 U590 ( .A(n508), .Z(n581) );
  NOR2_X1 U591 ( .A1(n578), .A2(n581), .ZN(n502) );
  XNOR2_X1 U592 ( .A(n502), .B(KEYINPUT104), .ZN(n503) );
  XNOR2_X1 U593 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n504) );
  XNOR2_X1 U594 ( .A(n565), .B(G119), .ZN(G21) );
  XNOR2_X1 U595 ( .A(KEYINPUT100), .B(n505), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n506) );
  XNOR2_X2 U597 ( .A(n506), .B(KEYINPUT102), .ZN(n589) );
  INV_X1 U598 ( .A(KEYINPUT106), .ZN(n507) );
  NOR2_X1 U599 ( .A1(n509), .A2(n508), .ZN(n510) );
  AND2_X1 U600 ( .A1(n591), .A2(n519), .ZN(n604) );
  AND2_X1 U601 ( .A1(n663), .A2(n512), .ZN(n513) );
  NAND2_X1 U602 ( .A1(n513), .A2(n578), .ZN(n514) );
  XNOR2_X1 U603 ( .A(n514), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U604 ( .A(n516), .B(n515), .ZN(n518) );
  NAND2_X1 U605 ( .A1(n518), .A2(n517), .ZN(n627) );
  XNOR2_X1 U606 ( .A(n627), .B(G140), .ZN(G42) );
  INV_X1 U607 ( .A(KEYINPUT53), .ZN(n638) );
  INV_X1 U608 ( .A(n525), .ZN(n527) );
  NAND2_X1 U609 ( .A1(n519), .A2(n527), .ZN(n520) );
  XNOR2_X1 U610 ( .A(n523), .B(KEYINPUT38), .ZN(n585) );
  INV_X1 U611 ( .A(n585), .ZN(n543) );
  NOR2_X2 U612 ( .A1(n543), .A2(n542), .ZN(n541) );
  NAND2_X1 U613 ( .A1(n541), .A2(n389), .ZN(n524) );
  NAND2_X1 U614 ( .A1(n563), .A2(n537), .ZN(n556) );
  OR2_X1 U615 ( .A1(n560), .A2(n525), .ZN(n526) );
  INV_X1 U616 ( .A(n560), .ZN(n592) );
  INV_X1 U617 ( .A(n578), .ZN(n608) );
  NOR2_X1 U618 ( .A1(n527), .A2(n608), .ZN(n528) );
  XOR2_X1 U619 ( .A(KEYINPUT50), .B(n528), .Z(n533) );
  NOR2_X1 U620 ( .A1(n529), .A2(n581), .ZN(n530) );
  XOR2_X1 U621 ( .A(KEYINPUT119), .B(n530), .Z(n531) );
  XNOR2_X1 U622 ( .A(KEYINPUT49), .B(n531), .ZN(n532) );
  NAND2_X1 U623 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U624 ( .A1(n592), .A2(n534), .ZN(n535) );
  NOR2_X1 U625 ( .A1(n348), .A2(n535), .ZN(n536) );
  XNOR2_X1 U626 ( .A(n536), .B(KEYINPUT51), .ZN(n538) );
  NAND2_X1 U627 ( .A1(n538), .A2(n537), .ZN(n550) );
  NOR2_X1 U628 ( .A1(n540), .A2(n539), .ZN(n677) );
  INV_X1 U629 ( .A(n677), .ZN(n625) );
  NAND2_X1 U630 ( .A1(n589), .A2(n625), .ZN(n614) );
  NAND2_X1 U631 ( .A1(n614), .A2(n541), .ZN(n547) );
  NAND2_X1 U632 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U633 ( .A(KEYINPUT120), .B(n544), .ZN(n545) );
  NAND2_X1 U634 ( .A1(n545), .A2(n389), .ZN(n546) );
  NAND2_X1 U635 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U636 ( .A1(n548), .A2(n563), .ZN(n549) );
  NAND2_X1 U637 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U638 ( .A(KEYINPUT52), .B(n551), .Z(n552) );
  NOR2_X1 U639 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U640 ( .A1(n554), .A2(G952), .ZN(n555) );
  NAND2_X1 U641 ( .A1(n556), .A2(n555), .ZN(n634) );
  XNOR2_X1 U642 ( .A(n557), .B(KEYINPUT22), .ZN(n558) );
  NAND2_X1 U643 ( .A1(n558), .A2(n578), .ZN(n559) );
  XNOR2_X1 U644 ( .A(n559), .B(KEYINPUT105), .ZN(n561) );
  NAND2_X1 U645 ( .A1(n561), .A2(n560), .ZN(n562) );
  INV_X1 U646 ( .A(n571), .ZN(n568) );
  NAND2_X1 U647 ( .A1(n565), .A2(n639), .ZN(n566) );
  INV_X1 U648 ( .A(KEYINPUT44), .ZN(n567) );
  NAND2_X1 U649 ( .A1(n348), .A2(n568), .ZN(n569) );
  OR2_X1 U650 ( .A1(n570), .A2(n592), .ZN(n572) );
  NOR2_X1 U651 ( .A1(n678), .A2(n345), .ZN(n573) );
  XNOR2_X1 U652 ( .A(n573), .B(KEYINPUT96), .ZN(n575) );
  INV_X1 U653 ( .A(n614), .ZN(n574) );
  XNOR2_X1 U654 ( .A(n576), .B(KEYINPUT103), .ZN(n583) );
  XNOR2_X1 U655 ( .A(n577), .B(KEYINPUT84), .ZN(n579) );
  NAND2_X1 U656 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U657 ( .A(n580), .B(KEYINPUT85), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n582), .A2(n581), .ZN(n662) );
  XNOR2_X1 U659 ( .A(KEYINPUT83), .B(KEYINPUT45), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n586), .A2(n585), .ZN(n588) );
  XNOR2_X1 U661 ( .A(n590), .B(KEYINPUT40), .ZN(n729) );
  INV_X1 U662 ( .A(n729), .ZN(n602) );
  XNOR2_X1 U663 ( .A(KEYINPUT28), .B(KEYINPUT111), .ZN(n594) );
  XNOR2_X1 U664 ( .A(n594), .B(n593), .ZN(n597) );
  XNOR2_X1 U665 ( .A(KEYINPUT110), .B(n595), .ZN(n596) );
  NOR2_X2 U666 ( .A1(n597), .A2(n596), .ZN(n612) );
  NAND2_X1 U667 ( .A1(n598), .A2(n612), .ZN(n600) );
  XOR2_X1 U668 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n599) );
  INV_X1 U669 ( .A(n726), .ZN(n601) );
  AND2_X1 U670 ( .A1(n604), .A2(n346), .ZN(n605) );
  NAND2_X1 U671 ( .A1(n663), .A2(n605), .ZN(n607) );
  XOR2_X1 U672 ( .A(KEYINPUT36), .B(KEYINPUT86), .Z(n606) );
  XNOR2_X1 U673 ( .A(n607), .B(n606), .ZN(n609) );
  NAND2_X1 U674 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U675 ( .A(n610), .B(KEYINPUT113), .ZN(n727) );
  NOR2_X1 U676 ( .A1(n611), .A2(n727), .ZN(n622) );
  NAND2_X1 U677 ( .A1(n672), .A2(n614), .ZN(n615) );
  OR2_X1 U678 ( .A1(KEYINPUT47), .A2(n615), .ZN(n620) );
  NAND2_X1 U679 ( .A1(n615), .A2(KEYINPUT47), .ZN(n617) );
  NAND2_X1 U680 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U681 ( .A(n618), .B(KEYINPUT81), .ZN(n619) );
  AND2_X1 U682 ( .A1(n620), .A2(n619), .ZN(n621) );
  AND2_X1 U683 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U684 ( .A(n623), .B(KEYINPUT48), .ZN(n629) );
  OR2_X1 U685 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U686 ( .A(n626), .B(KEYINPUT114), .ZN(n731) );
  AND2_X1 U687 ( .A1(n627), .A2(n731), .ZN(n628) );
  NAND2_X1 U688 ( .A1(n629), .A2(n628), .ZN(n718) );
  INV_X1 U689 ( .A(n718), .ZN(n630) );
  NOR2_X1 U690 ( .A1(n642), .A2(KEYINPUT2), .ZN(n631) );
  NOR2_X1 U691 ( .A1(n647), .A2(n631), .ZN(n632) );
  XNOR2_X1 U692 ( .A(n632), .B(KEYINPUT82), .ZN(n633) );
  NAND2_X1 U693 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U694 ( .A(n638), .B(n637), .ZN(G75) );
  XNOR2_X1 U695 ( .A(n639), .B(G122), .ZN(G24) );
  XOR2_X1 U696 ( .A(n640), .B(G110), .Z(G12) );
  AND2_X1 U697 ( .A1(KEYINPUT68), .A2(KEYINPUT2), .ZN(n641) );
  INV_X1 U698 ( .A(KEYINPUT2), .ZN(n643) );
  NOR2_X1 U699 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U700 ( .A1(n645), .A2(KEYINPUT68), .ZN(n646) );
  NAND2_X1 U701 ( .A1(n693), .A2(G472), .ZN(n650) );
  XNOR2_X1 U702 ( .A(n648), .B(KEYINPUT62), .ZN(n649) );
  XNOR2_X1 U703 ( .A(n650), .B(n649), .ZN(n651) );
  NAND2_X1 U704 ( .A1(n651), .A2(n659), .ZN(n654) );
  XNOR2_X1 U705 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n652) );
  XNOR2_X1 U706 ( .A(n652), .B(KEYINPUT87), .ZN(n653) );
  XNOR2_X1 U707 ( .A(n654), .B(n653), .ZN(G57) );
  NAND2_X1 U708 ( .A1(n693), .A2(G469), .ZN(n658) );
  XNOR2_X1 U709 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n655) );
  XNOR2_X1 U710 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U711 ( .A(n658), .B(n657), .ZN(n660) );
  INV_X1 U712 ( .A(n659), .ZN(n702) );
  NOR2_X2 U713 ( .A1(n660), .A2(n702), .ZN(n661) );
  XNOR2_X1 U714 ( .A(n661), .B(KEYINPUT122), .ZN(G54) );
  XNOR2_X1 U715 ( .A(G101), .B(n662), .ZN(G3) );
  NAND2_X1 U716 ( .A1(n345), .A2(n663), .ZN(n664) );
  XNOR2_X1 U717 ( .A(n664), .B(G104), .ZN(G6) );
  XOR2_X1 U718 ( .A(KEYINPUT27), .B(KEYINPUT116), .Z(n666) );
  XNOR2_X1 U719 ( .A(G107), .B(KEYINPUT26), .ZN(n665) );
  XNOR2_X1 U720 ( .A(n666), .B(n665), .ZN(n667) );
  XOR2_X1 U721 ( .A(KEYINPUT115), .B(n667), .Z(n669) );
  NAND2_X1 U722 ( .A1(n345), .A2(n677), .ZN(n668) );
  XNOR2_X1 U723 ( .A(n669), .B(n668), .ZN(G9) );
  XOR2_X1 U724 ( .A(G128), .B(KEYINPUT29), .Z(n671) );
  NAND2_X1 U725 ( .A1(n672), .A2(n677), .ZN(n670) );
  XNOR2_X1 U726 ( .A(n671), .B(n670), .ZN(G30) );
  XOR2_X1 U727 ( .A(G146), .B(KEYINPUT117), .Z(n674) );
  NAND2_X1 U728 ( .A1(n672), .A2(n663), .ZN(n673) );
  XNOR2_X1 U729 ( .A(n674), .B(n673), .ZN(G48) );
  NAND2_X1 U730 ( .A1(n678), .A2(n663), .ZN(n675) );
  XNOR2_X1 U731 ( .A(n675), .B(KEYINPUT118), .ZN(n676) );
  XNOR2_X1 U732 ( .A(G113), .B(n676), .ZN(G15) );
  NAND2_X1 U733 ( .A1(n678), .A2(n677), .ZN(n679) );
  XNOR2_X1 U734 ( .A(n679), .B(G116), .ZN(G18) );
  NAND2_X1 U735 ( .A1(n693), .A2(G210), .ZN(n685) );
  XOR2_X1 U736 ( .A(KEYINPUT54), .B(KEYINPUT121), .Z(n682) );
  XNOR2_X1 U737 ( .A(KEYINPUT88), .B(KEYINPUT55), .ZN(n681) );
  XNOR2_X1 U738 ( .A(n682), .B(n681), .ZN(n683) );
  XNOR2_X1 U739 ( .A(n680), .B(n683), .ZN(n684) );
  XNOR2_X1 U740 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X2 U741 ( .A1(n686), .A2(n702), .ZN(n687) );
  XNOR2_X1 U742 ( .A(n687), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U743 ( .A1(n693), .A2(G475), .ZN(n690) );
  XOR2_X1 U744 ( .A(n688), .B(KEYINPUT59), .Z(n689) );
  XNOR2_X1 U745 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X2 U746 ( .A1(n691), .A2(n702), .ZN(n692) );
  XNOR2_X1 U747 ( .A(n692), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U748 ( .A1(n697), .A2(G478), .ZN(n695) );
  XNOR2_X1 U749 ( .A(n695), .B(n694), .ZN(n696) );
  NOR2_X1 U750 ( .A1(n702), .A2(n696), .ZN(G63) );
  NAND2_X1 U751 ( .A1(n697), .A2(G217), .ZN(n700) );
  XOR2_X1 U752 ( .A(n698), .B(KEYINPUT123), .Z(n699) );
  XNOR2_X1 U753 ( .A(n700), .B(n699), .ZN(n701) );
  NOR2_X1 U754 ( .A1(n702), .A2(n701), .ZN(G66) );
  NOR2_X1 U755 ( .A1(n703), .A2(G953), .ZN(n708) );
  NAND2_X1 U756 ( .A1(G953), .A2(G224), .ZN(n704) );
  XNOR2_X1 U757 ( .A(KEYINPUT61), .B(n704), .ZN(n705) );
  NAND2_X1 U758 ( .A1(n705), .A2(G898), .ZN(n706) );
  XOR2_X1 U759 ( .A(KEYINPUT124), .B(n706), .Z(n707) );
  NOR2_X1 U760 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U761 ( .A(n709), .B(KEYINPUT125), .ZN(n714) );
  XOR2_X1 U762 ( .A(G101), .B(n710), .Z(n712) );
  NOR2_X1 U763 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U764 ( .A(n714), .B(n713), .ZN(G69) );
  XOR2_X1 U765 ( .A(n716), .B(n715), .Z(n717) );
  XNOR2_X1 U766 ( .A(KEYINPUT126), .B(n717), .ZN(n721) );
  XNOR2_X1 U767 ( .A(n721), .B(n718), .ZN(n720) );
  NAND2_X1 U768 ( .A1(n720), .A2(n719), .ZN(n725) );
  XNOR2_X1 U769 ( .A(G227), .B(n721), .ZN(n722) );
  NAND2_X1 U770 ( .A1(n722), .A2(G900), .ZN(n723) );
  NAND2_X1 U771 ( .A1(G953), .A2(n723), .ZN(n724) );
  NAND2_X1 U772 ( .A1(n725), .A2(n724), .ZN(G72) );
  XOR2_X1 U773 ( .A(n726), .B(G137), .Z(G39) );
  XNOR2_X1 U774 ( .A(n727), .B(G125), .ZN(n728) );
  XNOR2_X1 U775 ( .A(n728), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U776 ( .A(G131), .B(KEYINPUT127), .ZN(n730) );
  XNOR2_X1 U777 ( .A(n730), .B(n729), .ZN(G33) );
  XNOR2_X1 U778 ( .A(G134), .B(n731), .ZN(G36) );
endmodule

