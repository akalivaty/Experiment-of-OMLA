

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U322 ( .A(n438), .B(n437), .ZN(n440) );
  XOR2_X1 U323 ( .A(KEYINPUT38), .B(n467), .Z(n494) );
  XOR2_X1 U324 ( .A(KEYINPUT28), .B(n458), .Z(n529) );
  XOR2_X1 U325 ( .A(G169GAT), .B(G176GAT), .Z(n290) );
  XOR2_X1 U326 ( .A(n434), .B(n433), .Z(n291) );
  NOR2_X1 U327 ( .A1(n400), .A2(n399), .ZN(n401) );
  XNOR2_X1 U328 ( .A(n436), .B(n290), .ZN(n437) );
  XNOR2_X1 U329 ( .A(KEYINPUT118), .B(KEYINPUT54), .ZN(n409) );
  XNOR2_X1 U330 ( .A(n354), .B(n365), .ZN(n355) );
  XNOR2_X1 U331 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U332 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U333 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n359) );
  XNOR2_X1 U334 ( .A(n573), .B(n359), .ZN(n544) );
  INV_X1 U335 ( .A(G43GAT), .ZN(n468) );
  XNOR2_X1 U336 ( .A(n444), .B(n443), .ZN(n527) );
  XNOR2_X1 U337 ( .A(n447), .B(G183GAT), .ZN(n448) );
  XNOR2_X1 U338 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U339 ( .A(n449), .B(n448), .ZN(G1350GAT) );
  XNOR2_X1 U340 ( .A(n471), .B(n470), .ZN(G1330GAT) );
  XOR2_X1 U341 ( .A(G85GAT), .B(G148GAT), .Z(n293) );
  XNOR2_X1 U342 ( .A(G141GAT), .B(G162GAT), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U344 ( .A(KEYINPUT5), .B(KEYINPUT90), .Z(n295) );
  XNOR2_X1 U345 ( .A(G127GAT), .B(G120GAT), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U347 ( .A(n297), .B(n296), .Z(n302) );
  XOR2_X1 U348 ( .A(KEYINPUT89), .B(KEYINPUT1), .Z(n299) );
  NAND2_X1 U349 ( .A1(G225GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U351 ( .A(G1GAT), .B(n300), .ZN(n301) );
  XNOR2_X1 U352 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U353 ( .A(KEYINPUT88), .B(KEYINPUT6), .Z(n304) );
  XNOR2_X1 U354 ( .A(G57GAT), .B(KEYINPUT4), .ZN(n303) );
  XNOR2_X1 U355 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U356 ( .A(n306), .B(n305), .Z(n311) );
  XOR2_X1 U357 ( .A(KEYINPUT80), .B(KEYINPUT0), .Z(n308) );
  XNOR2_X1 U358 ( .A(G113GAT), .B(G134GAT), .ZN(n307) );
  XNOR2_X1 U359 ( .A(n308), .B(n307), .ZN(n436) );
  XNOR2_X1 U360 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n309), .B(KEYINPUT3), .ZN(n422) );
  XNOR2_X1 U362 ( .A(n436), .B(n422), .ZN(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n489) );
  XNOR2_X1 U364 ( .A(G29GAT), .B(n489), .ZN(n514) );
  XOR2_X1 U365 ( .A(G211GAT), .B(G218GAT), .Z(n313) );
  XNOR2_X1 U366 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U368 ( .A(G197GAT), .B(n314), .ZN(n428) );
  XOR2_X1 U369 ( .A(G183GAT), .B(KEYINPUT19), .Z(n316) );
  XNOR2_X1 U370 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n433) );
  XOR2_X1 U372 ( .A(n433), .B(KEYINPUT91), .Z(n318) );
  NAND2_X1 U373 ( .A1(G226GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U375 ( .A(G36GAT), .B(G190GAT), .Z(n394) );
  XOR2_X1 U376 ( .A(n319), .B(n394), .Z(n322) );
  XOR2_X1 U377 ( .A(G169GAT), .B(G8GAT), .Z(n329) );
  XNOR2_X1 U378 ( .A(G176GAT), .B(G92GAT), .ZN(n320) );
  XNOR2_X1 U379 ( .A(n320), .B(G64GAT), .ZN(n346) );
  XNOR2_X1 U380 ( .A(n329), .B(n346), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U382 ( .A(n428), .B(n323), .Z(n517) );
  XOR2_X1 U383 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n325) );
  XNOR2_X1 U384 ( .A(KEYINPUT71), .B(KEYINPUT70), .ZN(n324) );
  XNOR2_X1 U385 ( .A(n325), .B(n324), .ZN(n342) );
  XOR2_X1 U386 ( .A(G1GAT), .B(G113GAT), .Z(n327) );
  XNOR2_X1 U387 ( .A(G197GAT), .B(G15GAT), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U389 ( .A(n328), .B(G50GAT), .Z(n331) );
  XNOR2_X1 U390 ( .A(n329), .B(G36GAT), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U392 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n333) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U395 ( .A(n335), .B(n334), .Z(n340) );
  XOR2_X1 U396 ( .A(KEYINPUT8), .B(KEYINPUT69), .Z(n337) );
  XNOR2_X1 U397 ( .A(G43GAT), .B(G29GAT), .ZN(n336) );
  XNOR2_X1 U398 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U399 ( .A(KEYINPUT7), .B(n338), .Z(n398) );
  XOR2_X1 U400 ( .A(G141GAT), .B(G22GAT), .Z(n412) );
  XNOR2_X1 U401 ( .A(n398), .B(n412), .ZN(n339) );
  XNOR2_X1 U402 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U403 ( .A(n342), .B(n341), .ZN(n568) );
  INV_X1 U404 ( .A(n568), .ZN(n555) );
  XOR2_X1 U405 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n344) );
  XNOR2_X1 U406 ( .A(G204GAT), .B(KEYINPUT74), .ZN(n343) );
  XNOR2_X1 U407 ( .A(n344), .B(n343), .ZN(n358) );
  XNOR2_X1 U408 ( .A(G106GAT), .B(G78GAT), .ZN(n345) );
  XNOR2_X1 U409 ( .A(n345), .B(G148GAT), .ZN(n413) );
  XNOR2_X1 U410 ( .A(n413), .B(n346), .ZN(n352) );
  XOR2_X1 U411 ( .A(KEYINPUT32), .B(KEYINPUT75), .Z(n348) );
  NAND2_X1 U412 ( .A1(G230GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U413 ( .A(n348), .B(n347), .ZN(n350) );
  INV_X1 U414 ( .A(KEYINPUT73), .ZN(n349) );
  XNOR2_X1 U415 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U417 ( .A(G120GAT), .B(G71GAT), .Z(n434) );
  XOR2_X1 U418 ( .A(G99GAT), .B(G85GAT), .Z(n391) );
  XOR2_X1 U419 ( .A(n434), .B(n391), .Z(n354) );
  XNOR2_X1 U420 ( .A(G57GAT), .B(KEYINPUT72), .ZN(n353) );
  XNOR2_X1 U421 ( .A(n353), .B(KEYINPUT13), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n358), .B(n357), .ZN(n573) );
  INV_X1 U423 ( .A(n544), .ZN(n496) );
  NAND2_X1 U424 ( .A1(n555), .A2(n496), .ZN(n360) );
  NAND2_X1 U425 ( .A1(KEYINPUT46), .A2(n360), .ZN(n364) );
  INV_X1 U426 ( .A(KEYINPUT46), .ZN(n361) );
  NAND2_X1 U427 ( .A1(n496), .A2(n361), .ZN(n362) );
  OR2_X1 U428 ( .A1(n568), .A2(n362), .ZN(n363) );
  AND2_X1 U429 ( .A1(n364), .A2(n363), .ZN(n400) );
  XOR2_X1 U430 ( .A(G15GAT), .B(G127GAT), .Z(n439) );
  XOR2_X1 U431 ( .A(n365), .B(n439), .Z(n367) );
  NAND2_X1 U432 ( .A1(G231GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U433 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U434 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n369) );
  XNOR2_X1 U435 ( .A(G64GAT), .B(KEYINPUT15), .ZN(n368) );
  XNOR2_X1 U436 ( .A(n369), .B(n368), .ZN(n370) );
  XOR2_X1 U437 ( .A(n371), .B(n370), .Z(n379) );
  XOR2_X1 U438 ( .A(G78GAT), .B(G155GAT), .Z(n373) );
  XNOR2_X1 U439 ( .A(G22GAT), .B(G211GAT), .ZN(n372) );
  XNOR2_X1 U440 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U441 ( .A(G183GAT), .B(G71GAT), .Z(n375) );
  XNOR2_X1 U442 ( .A(G8GAT), .B(G1GAT), .ZN(n374) );
  XNOR2_X1 U443 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U444 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U445 ( .A(n379), .B(n378), .Z(n533) );
  INV_X1 U446 ( .A(n533), .ZN(n577) );
  XOR2_X1 U447 ( .A(G92GAT), .B(G106GAT), .Z(n381) );
  XNOR2_X1 U448 ( .A(G134GAT), .B(G218GAT), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U450 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n383) );
  XNOR2_X1 U451 ( .A(KEYINPUT78), .B(KEYINPUT9), .ZN(n382) );
  XNOR2_X1 U452 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U453 ( .A(n385), .B(n384), .Z(n390) );
  XOR2_X1 U454 ( .A(KEYINPUT66), .B(KEYINPUT77), .Z(n387) );
  NAND2_X1 U455 ( .A1(G232GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U456 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U457 ( .A(KEYINPUT65), .B(n388), .ZN(n389) );
  XNOR2_X1 U458 ( .A(n390), .B(n389), .ZN(n392) );
  XOR2_X1 U459 ( .A(n392), .B(n391), .Z(n396) );
  XNOR2_X1 U460 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n393) );
  XNOR2_X1 U461 ( .A(n393), .B(G162GAT), .ZN(n423) );
  XNOR2_X1 U462 ( .A(n423), .B(n394), .ZN(n395) );
  XNOR2_X1 U463 ( .A(n396), .B(n395), .ZN(n397) );
  XOR2_X1 U464 ( .A(n398), .B(n397), .Z(n553) );
  INV_X1 U465 ( .A(n553), .ZN(n561) );
  NAND2_X1 U466 ( .A1(n577), .A2(n553), .ZN(n399) );
  XNOR2_X1 U467 ( .A(n401), .B(KEYINPUT47), .ZN(n407) );
  XOR2_X1 U468 ( .A(KEYINPUT45), .B(KEYINPUT110), .Z(n403) );
  XOR2_X1 U469 ( .A(KEYINPUT36), .B(n561), .Z(n582) );
  NOR2_X1 U470 ( .A1(n577), .A2(n582), .ZN(n402) );
  XNOR2_X1 U471 ( .A(n403), .B(n402), .ZN(n404) );
  NOR2_X1 U472 ( .A1(n573), .A2(n404), .ZN(n405) );
  NAND2_X1 U473 ( .A1(n405), .A2(n568), .ZN(n406) );
  NAND2_X1 U474 ( .A1(n407), .A2(n406), .ZN(n408) );
  XNOR2_X1 U475 ( .A(n408), .B(KEYINPUT48), .ZN(n524) );
  NAND2_X1 U476 ( .A1(n517), .A2(n524), .ZN(n410) );
  NOR2_X1 U477 ( .A1(n514), .A2(n411), .ZN(n567) );
  XOR2_X1 U478 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U479 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U480 ( .A(n415), .B(n414), .ZN(n427) );
  XOR2_X1 U481 ( .A(KEYINPUT23), .B(KEYINPUT84), .Z(n417) );
  XNOR2_X1 U482 ( .A(KEYINPUT85), .B(KEYINPUT83), .ZN(n416) );
  XNOR2_X1 U483 ( .A(n417), .B(n416), .ZN(n421) );
  XOR2_X1 U484 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n419) );
  XNOR2_X1 U485 ( .A(KEYINPUT87), .B(KEYINPUT86), .ZN(n418) );
  XNOR2_X1 U486 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U487 ( .A(n421), .B(n420), .Z(n425) );
  XNOR2_X1 U488 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U489 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n429) );
  XNOR2_X1 U491 ( .A(n429), .B(n428), .ZN(n458) );
  NAND2_X1 U492 ( .A1(n567), .A2(n458), .ZN(n430) );
  XNOR2_X1 U493 ( .A(n430), .B(KEYINPUT55), .ZN(n445) );
  XOR2_X1 U494 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n432) );
  XNOR2_X1 U495 ( .A(G43GAT), .B(KEYINPUT20), .ZN(n431) );
  XNOR2_X1 U496 ( .A(n432), .B(n431), .ZN(n444) );
  NAND2_X1 U497 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U498 ( .A(n291), .B(n435), .ZN(n438) );
  XOR2_X1 U499 ( .A(n440), .B(n439), .Z(n442) );
  XNOR2_X1 U500 ( .A(G99GAT), .B(G190GAT), .ZN(n441) );
  XNOR2_X1 U501 ( .A(n442), .B(n441), .ZN(n443) );
  NAND2_X1 U502 ( .A1(n445), .A2(n527), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n446), .B(KEYINPUT119), .ZN(n562) );
  NAND2_X1 U504 ( .A1(n562), .A2(n533), .ZN(n449) );
  XOR2_X1 U505 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n447) );
  NOR2_X1 U506 ( .A1(n527), .A2(n458), .ZN(n450) );
  XNOR2_X1 U507 ( .A(KEYINPUT26), .B(n450), .ZN(n566) );
  XNOR2_X1 U508 ( .A(KEYINPUT27), .B(n517), .ZN(n459) );
  NAND2_X1 U509 ( .A1(n566), .A2(n459), .ZN(n451) );
  XNOR2_X1 U510 ( .A(n451), .B(KEYINPUT93), .ZN(n456) );
  NAND2_X1 U511 ( .A1(n527), .A2(n517), .ZN(n452) );
  NAND2_X1 U512 ( .A1(n452), .A2(n458), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n453), .B(KEYINPUT94), .ZN(n454) );
  XNOR2_X1 U514 ( .A(KEYINPUT25), .B(n454), .ZN(n455) );
  NOR2_X1 U515 ( .A1(n456), .A2(n455), .ZN(n457) );
  NOR2_X1 U516 ( .A1(n457), .A2(n514), .ZN(n464) );
  INV_X1 U517 ( .A(n529), .ZN(n461) );
  NAND2_X1 U518 ( .A1(n514), .A2(n459), .ZN(n460) );
  XOR2_X1 U519 ( .A(KEYINPUT92), .B(n460), .Z(n525) );
  NAND2_X1 U520 ( .A1(n461), .A2(n525), .ZN(n462) );
  NOR2_X1 U521 ( .A1(n462), .A2(n527), .ZN(n463) );
  NOR2_X1 U522 ( .A1(n464), .A2(n463), .ZN(n475) );
  NOR2_X1 U523 ( .A1(n582), .A2(n475), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n577), .A2(n465), .ZN(n466) );
  XNOR2_X1 U525 ( .A(KEYINPUT37), .B(n466), .ZN(n511) );
  NOR2_X1 U526 ( .A1(n568), .A2(n573), .ZN(n476) );
  NAND2_X1 U527 ( .A1(n511), .A2(n476), .ZN(n467) );
  NAND2_X1 U528 ( .A1(n494), .A2(n527), .ZN(n471) );
  XOR2_X1 U529 ( .A(KEYINPUT40), .B(KEYINPUT100), .Z(n469) );
  XOR2_X1 U530 ( .A(KEYINPUT96), .B(KEYINPUT34), .Z(n479) );
  XOR2_X1 U531 ( .A(KEYINPUT79), .B(KEYINPUT16), .Z(n473) );
  NAND2_X1 U532 ( .A1(n553), .A2(n533), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n473), .B(n472), .ZN(n474) );
  NOR2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n498) );
  NAND2_X1 U535 ( .A1(n498), .A2(n476), .ZN(n477) );
  XNOR2_X1 U536 ( .A(n477), .B(KEYINPUT95), .ZN(n486) );
  NAND2_X1 U537 ( .A1(n486), .A2(n514), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U539 ( .A(G1GAT), .B(n480), .Z(G1324GAT) );
  XOR2_X1 U540 ( .A(G8GAT), .B(KEYINPUT97), .Z(n482) );
  NAND2_X1 U541 ( .A1(n486), .A2(n517), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT98), .B(KEYINPUT35), .Z(n484) );
  NAND2_X1 U544 ( .A1(n486), .A2(n527), .ZN(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(n485), .ZN(G1326GAT) );
  XOR2_X1 U547 ( .A(G22GAT), .B(KEYINPUT99), .Z(n488) );
  NAND2_X1 U548 ( .A1(n486), .A2(n529), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(G1327GAT) );
  NAND2_X1 U550 ( .A1(n489), .A2(n494), .ZN(n491) );
  OR2_X1 U551 ( .A1(n494), .A2(G29GAT), .ZN(n490) );
  NAND2_X1 U552 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U553 ( .A(KEYINPUT39), .B(n492), .ZN(G1328GAT) );
  NAND2_X1 U554 ( .A1(n494), .A2(n517), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n493), .B(G36GAT), .ZN(G1329GAT) );
  AND2_X1 U556 ( .A1(n529), .A2(n494), .ZN(n495) );
  XOR2_X1 U557 ( .A(G50GAT), .B(n495), .Z(G1331GAT) );
  NAND2_X1 U558 ( .A1(n568), .A2(n496), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n497), .B(KEYINPUT101), .ZN(n512) );
  AND2_X1 U560 ( .A1(n512), .A2(n498), .ZN(n508) );
  NAND2_X1 U561 ( .A1(n514), .A2(n508), .ZN(n501) );
  XNOR2_X1 U562 ( .A(G57GAT), .B(KEYINPUT102), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(KEYINPUT42), .ZN(n500) );
  XNOR2_X1 U564 ( .A(n501), .B(n500), .ZN(G1332GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n503) );
  NAND2_X1 U566 ( .A1(n508), .A2(n517), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G64GAT), .B(n504), .ZN(G1333GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n506) );
  NAND2_X1 U570 ( .A1(n508), .A2(n527), .ZN(n505) );
  XNOR2_X1 U571 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U572 ( .A(G71GAT), .B(n507), .ZN(G1334GAT) );
  XOR2_X1 U573 ( .A(G78GAT), .B(KEYINPUT43), .Z(n510) );
  NAND2_X1 U574 ( .A1(n508), .A2(n529), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NAND2_X1 U576 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(KEYINPUT107), .ZN(n521) );
  NAND2_X1 U578 ( .A1(n514), .A2(n521), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n515), .B(KEYINPUT108), .ZN(n516) );
  XNOR2_X1 U580 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n517), .A2(n521), .ZN(n518) );
  XNOR2_X1 U582 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U583 ( .A(G99GAT), .B(KEYINPUT109), .Z(n520) );
  NAND2_X1 U584 ( .A1(n521), .A2(n527), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n520), .B(n519), .ZN(G1338GAT) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n523) );
  NAND2_X1 U587 ( .A1(n521), .A2(n529), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(G1339GAT) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(KEYINPUT111), .ZN(n541) );
  NAND2_X1 U591 ( .A1(n541), .A2(n527), .ZN(n528) );
  NOR2_X1 U592 ( .A1(n529), .A2(n528), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n555), .A2(n537), .ZN(n530) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(G120GAT), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U596 ( .A1(n537), .A2(n496), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT112), .B(KEYINPUT50), .Z(n535) );
  NAND2_X1 U599 ( .A1(n537), .A2(n533), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U601 ( .A(G127GAT), .B(n536), .Z(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U603 ( .A1(n537), .A2(n561), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U605 ( .A(G134GAT), .B(n540), .Z(G1343GAT) );
  NAND2_X1 U606 ( .A1(n541), .A2(n566), .ZN(n552) );
  NOR2_X1 U607 ( .A1(n568), .A2(n552), .ZN(n542) );
  XOR2_X1 U608 ( .A(G141GAT), .B(n542), .Z(n543) );
  XNOR2_X1 U609 ( .A(KEYINPUT114), .B(n543), .ZN(G1344GAT) );
  NOR2_X1 U610 ( .A1(n544), .A2(n552), .ZN(n549) );
  XOR2_X1 U611 ( .A(KEYINPUT116), .B(KEYINPUT53), .Z(n546) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(KEYINPUT115), .B(n547), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n549), .B(n548), .ZN(G1345GAT) );
  NOR2_X1 U616 ( .A1(n577), .A2(n552), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(KEYINPUT117), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1346GAT) );
  NOR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U620 ( .A(G162GAT), .B(n554), .Z(G1347GAT) );
  NAND2_X1 U621 ( .A1(n562), .A2(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n556), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n562), .A2(n496), .ZN(n558) );
  XOR2_X1 U624 ( .A(KEYINPUT120), .B(KEYINPUT57), .Z(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1349GAT) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT58), .B(KEYINPUT123), .Z(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n565), .B(G190GAT), .ZN(G1351GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n581) );
  NOR2_X1 U633 ( .A1(n568), .A2(n581), .ZN(n572) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT60), .B(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  INV_X1 U638 ( .A(n573), .ZN(n574) );
  NOR2_X1 U639 ( .A1(n574), .A2(n581), .ZN(n576) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n581), .ZN(n578) );
  XOR2_X1 U643 ( .A(G211GAT), .B(n578), .Z(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT125), .B(KEYINPUT62), .Z(n580) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n579) );
  XNOR2_X1 U646 ( .A(n580), .B(n579), .ZN(n584) );
  NOR2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U648 ( .A(n584), .B(n583), .Z(G1355GAT) );
endmodule

