//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 0 0 1 0 1 1 0 1 0 1 1 0 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0 0 1 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:16 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n636, new_n638, new_n639, new_n640,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g019(.A(KEYINPUT65), .B(G452), .ZN(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT66), .Z(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n452), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(G2106), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT67), .Z(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT68), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G125), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n462), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n464), .A2(new_n466), .A3(G137), .ZN(new_n475));
  NAND2_X1  g050(.A1(G101), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT69), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NOR3_X1   g054(.A1(new_n474), .A2(KEYINPUT69), .A3(new_n477), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n467), .A2(new_n462), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n467), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  AND3_X1   g064(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT68), .ZN(new_n490));
  AOI21_X1  g065(.A(KEYINPUT68), .B1(new_n464), .B2(new_n466), .ZN(new_n491));
  OAI211_X1 g066(.A(G138), .B(new_n462), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n464), .A2(new_n466), .A3(KEYINPUT4), .A4(G138), .ZN(new_n495));
  NAND2_X1  g070(.A1(G102), .A2(G2104), .ZN(new_n496));
  AOI21_X1  g071(.A(G2105), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n464), .A2(new_n466), .A3(G126), .ZN(new_n498));
  NAND2_X1  g073(.A1(G114), .A2(G2104), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n462), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n494), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI211_X1 g087(.A(new_n508), .B(new_n510), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n505), .A2(new_n506), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n508), .A2(new_n510), .ZN(new_n516));
  INV_X1    g091(.A(G62), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT70), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(G75), .A2(G543), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT5), .B(G543), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(new_n521), .A3(G62), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n518), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n515), .B1(new_n523), .B2(G651), .ZN(G166));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  INV_X1    g100(.A(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT71), .B(G89), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  OAI221_X1 g104(.A(new_n527), .B1(new_n513), .B2(new_n528), .C1(new_n505), .C2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n520), .A2(G63), .ZN(new_n532));
  NAND3_X1  g107(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n530), .A2(new_n534), .ZN(G168));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  INV_X1    g111(.A(G64), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n536), .B1(new_n516), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G651), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(G52), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  OAI22_X1  g118(.A1(new_n505), .A2(new_n542), .B1(new_n513), .B2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n538), .A2(KEYINPUT72), .A3(G651), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n541), .A2(new_n545), .A3(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  AOI22_X1  g123(.A1(new_n520), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n549), .A2(new_n531), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n504), .A2(G43), .A3(G543), .ZN(new_n551));
  INV_X1    g126(.A(G81), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n552), .B2(new_n513), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT73), .Z(G188));
  OAI211_X1 g136(.A(G53), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n562));
  OR2_X1    g137(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(KEYINPUT74), .A2(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G91), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n566), .A2(new_n513), .B1(new_n562), .B2(new_n564), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(KEYINPUT75), .ZN(new_n570));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G65), .ZN(new_n572));
  NAND4_X1  g147(.A1(new_n508), .A2(new_n510), .A3(new_n570), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(G78), .A2(G543), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g150(.A(KEYINPUT76), .B1(new_n575), .B2(G651), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  AOI211_X1 g152(.A(new_n577), .B(new_n531), .C1(new_n573), .C2(new_n574), .ZN(new_n578));
  OAI211_X1 g153(.A(new_n565), .B(new_n568), .C1(new_n576), .C2(new_n578), .ZN(G299));
  NAND2_X1  g154(.A1(new_n532), .A2(new_n533), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(G651), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n504), .A2(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G51), .ZN(new_n583));
  OR2_X1    g158(.A1(new_n513), .A2(new_n528), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n581), .A2(new_n583), .A3(new_n527), .A4(new_n584), .ZN(G286));
  NAND2_X1  g160(.A1(new_n523), .A2(G651), .ZN(new_n586));
  INV_X1    g161(.A(new_n515), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G303));
  OAI21_X1  g163(.A(G651), .B1(new_n520), .B2(G74), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT77), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n520), .A2(new_n504), .A3(G87), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n504), .A2(G49), .A3(G543), .ZN(new_n593));
  OAI211_X1 g168(.A(KEYINPUT77), .B(G651), .C1(new_n520), .C2(G74), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n591), .A2(new_n592), .A3(new_n593), .A4(new_n594), .ZN(G288));
  INV_X1    g170(.A(G48), .ZN(new_n596));
  INV_X1    g171(.A(G86), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n505), .A2(new_n596), .B1(new_n513), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(G73), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G61), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n516), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n602), .A2(KEYINPUT78), .A3(G651), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  AOI21_X1  g179(.A(KEYINPUT78), .B1(new_n602), .B2(G651), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n599), .B1(new_n604), .B2(new_n605), .ZN(G305));
  AOI22_X1  g181(.A1(new_n520), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(new_n531), .ZN(new_n608));
  INV_X1    g183(.A(G47), .ZN(new_n609));
  INV_X1    g184(.A(G85), .ZN(new_n610));
  OAI22_X1  g185(.A1(new_n505), .A2(new_n609), .B1(new_n513), .B2(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  INV_X1    g190(.A(G66), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n516), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G651), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n582), .A2(G54), .ZN(new_n619));
  INV_X1    g194(.A(G92), .ZN(new_n620));
  OAI21_X1  g195(.A(KEYINPUT10), .B1(new_n513), .B2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n622));
  NAND4_X1  g197(.A1(new_n520), .A2(new_n504), .A3(new_n622), .A4(G92), .ZN(new_n623));
  AND4_X1   g198(.A1(new_n618), .A2(new_n619), .A3(new_n621), .A4(new_n623), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n614), .B1(G868), .B2(new_n624), .ZN(G284));
  OAI21_X1  g200(.A(new_n614), .B1(G868), .B2(new_n624), .ZN(G321));
  NAND2_X1  g201(.A1(G286), .A2(G868), .ZN(new_n627));
  INV_X1    g202(.A(new_n565), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT75), .B(G65), .ZN(new_n629));
  AOI22_X1  g204(.A1(new_n520), .A2(new_n629), .B1(G78), .B2(G543), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n577), .B1(new_n630), .B2(new_n531), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n575), .A2(KEYINPUT76), .A3(G651), .ZN(new_n632));
  AOI211_X1 g207(.A(new_n567), .B(new_n628), .C1(new_n631), .C2(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n627), .B1(new_n633), .B2(G868), .ZN(G297));
  OAI21_X1  g209(.A(new_n627), .B1(new_n633), .B2(G868), .ZN(G280));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n624), .B1(new_n636), .B2(G860), .ZN(G148));
  NAND2_X1  g212(.A1(new_n624), .A2(new_n636), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT79), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(G868), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n640), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g216(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g217(.A1(new_n471), .A2(G2104), .A3(new_n462), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT12), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT13), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2100), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n462), .A2(G111), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT80), .Z(new_n648));
  OAI211_X1 g223(.A(new_n648), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n484), .A2(G135), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n482), .A2(G123), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(G2096), .Z(new_n653));
  NAND2_X1  g228(.A1(new_n646), .A2(new_n653), .ZN(G156));
  XNOR2_X1  g229(.A(KEYINPUT15), .B(G2435), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT82), .B(G2438), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(G2427), .B(G2430), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT14), .ZN(new_n660));
  XOR2_X1   g235(.A(KEYINPUT81), .B(KEYINPUT16), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(G2451), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(G2454), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2443), .B(G2446), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n666), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1341), .B(G1348), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n667), .A2(new_n670), .A3(new_n668), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n672), .A2(G14), .A3(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(G401));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  XOR2_X1   g251(.A(G2067), .B(G2678), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G2084), .B(G2090), .Z(new_n679));
  NAND2_X1  g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n676), .B1(new_n680), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G2096), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n678), .A2(new_n679), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n686), .A2(new_n680), .A3(KEYINPUT17), .ZN(new_n687));
  AND2_X1   g262(.A1(new_n687), .A2(new_n681), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n685), .B(new_n688), .Z(G227));
  XNOR2_X1  g264(.A(KEYINPUT22), .B(G1981), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(G1971), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT19), .ZN(new_n693));
  XOR2_X1   g268(.A(G1956), .B(G2474), .Z(new_n694));
  XOR2_X1   g269(.A(G1961), .B(G1966), .Z(new_n695));
  NAND2_X1  g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT85), .ZN(new_n698));
  INV_X1    g273(.A(KEYINPUT84), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n698), .A2(new_n699), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT20), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n694), .A2(new_n695), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(new_n696), .ZN(new_n706));
  MUX2_X1   g281(.A(new_n705), .B(new_n706), .S(new_n693), .Z(new_n707));
  NAND3_X1  g282(.A1(new_n700), .A2(new_n701), .A3(KEYINPUT20), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n704), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT21), .B(G1986), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n704), .A2(new_n707), .A3(new_n708), .A4(new_n710), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n714), .B1(new_n712), .B2(new_n715), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n691), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n712), .A2(new_n715), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(new_n713), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n721), .A2(new_n690), .A3(new_n716), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n719), .A2(new_n722), .ZN(G229));
  AOI22_X1  g298(.A1(G119), .A2(new_n482), .B1(new_n484), .B2(G131), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n725));
  NOR2_X1   g300(.A1(G95), .A2(G2105), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT86), .Z(new_n727));
  OAI21_X1  g302(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G25), .B(new_n728), .S(G29), .Z(new_n729));
  XNOR2_X1  g304(.A(KEYINPUT35), .B(G1991), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n729), .B(new_n730), .Z(new_n731));
  INV_X1    g306(.A(G16), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G24), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n733), .B1(new_n612), .B2(new_n732), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT87), .B(G1986), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n734), .B(new_n735), .Z(new_n736));
  INV_X1    g311(.A(KEYINPUT91), .ZN(new_n737));
  INV_X1    g312(.A(KEYINPUT36), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n731), .B(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  INV_X1    g314(.A(KEYINPUT34), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n732), .A2(G23), .ZN(new_n741));
  INV_X1    g316(.A(G288), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n741), .B1(new_n742), .B2(new_n732), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT88), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT33), .B(G1976), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(KEYINPUT88), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n743), .B(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(new_n745), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n746), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n732), .A2(G6), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n602), .A2(G651), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT78), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n598), .B1(new_n755), .B2(new_n603), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n752), .B1(new_n756), .B2(new_n732), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT32), .B(G1981), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n732), .A2(G22), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G166), .B2(new_n732), .ZN(new_n761));
  XOR2_X1   g336(.A(KEYINPUT89), .B(G1971), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT90), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n761), .B(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n740), .B1(new_n751), .B2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n765), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n767), .A2(KEYINPUT34), .A3(new_n746), .A4(new_n750), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n739), .B1(new_n766), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n737), .A2(new_n738), .ZN(new_n770));
  NOR2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n624), .A2(G16), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G4), .B2(G16), .ZN(new_n773));
  INV_X1    g348(.A(G1348), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  INV_X1    g351(.A(KEYINPUT24), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n777), .A2(G34), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n777), .A2(G34), .ZN(new_n780));
  AOI21_X1  g355(.A(G29), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G29), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(G160), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n776), .B1(new_n784), .B2(G2084), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n732), .A2(G5), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(G171), .B2(new_n732), .ZN(new_n787));
  INV_X1    g362(.A(G1961), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  OR3_X1    g364(.A1(new_n474), .A2(KEYINPUT69), .A3(new_n477), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(new_n478), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n781), .B1(new_n791), .B2(G29), .ZN(new_n792));
  INV_X1    g367(.A(G2084), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n488), .A2(G29), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT29), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n783), .A2(G35), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n795), .B1(new_n794), .B2(new_n796), .ZN(new_n798));
  OR3_X1    g373(.A1(new_n797), .A2(new_n798), .A3(G2090), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT99), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n792), .A2(new_n793), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AND4_X1   g376(.A1(new_n775), .A2(new_n785), .A3(new_n789), .A4(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n652), .A2(new_n783), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT97), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n732), .A2(G19), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n554), .B2(new_n732), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1341), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n773), .A2(new_n774), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT30), .B(G28), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n809), .B1(new_n783), .B2(new_n810), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n808), .B(new_n811), .C1(new_n800), .C2(new_n799), .ZN(new_n812));
  INV_X1    g387(.A(G27), .ZN(new_n813));
  OAI21_X1  g388(.A(KEYINPUT98), .B1(new_n813), .B2(G29), .ZN(new_n814));
  OR3_X1    g389(.A1(new_n813), .A2(KEYINPUT98), .A3(G29), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n814), .B(new_n815), .C1(G164), .C2(new_n783), .ZN(new_n816));
  INV_X1    g391(.A(G2078), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n484), .A2(G139), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT25), .Z(new_n821));
  AOI22_X1  g396(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n819), .B(new_n821), .C1(new_n822), .C2(new_n462), .ZN(new_n823));
  MUX2_X1   g398(.A(G33), .B(new_n823), .S(G29), .Z(new_n824));
  NAND2_X1  g399(.A1(G168), .A2(G16), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n825), .B1(G16), .B2(G21), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT95), .B(G1966), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n824), .A2(G2072), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n818), .B(new_n829), .C1(G2072), .C2(new_n824), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n812), .A2(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n832));
  OAI21_X1  g407(.A(G2090), .B1(new_n797), .B2(new_n798), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT100), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n732), .A2(KEYINPUT23), .A3(G20), .ZN(new_n836));
  AOI21_X1  g411(.A(KEYINPUT23), .B1(new_n732), .B2(G20), .ZN(new_n837));
  AOI211_X1 g412(.A(new_n836), .B(new_n837), .C1(G299), .C2(G16), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G1956), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n832), .B1(new_n835), .B2(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n835), .A2(new_n832), .A3(new_n839), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n802), .B(new_n831), .C1(new_n840), .C2(new_n842), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n771), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n484), .A2(G141), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT92), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n848));
  NAND3_X1  g423(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT26), .ZN(new_n850));
  AOI211_X1 g425(.A(new_n848), .B(new_n850), .C1(G129), .C2(new_n482), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n847), .A2(G29), .A3(new_n851), .ZN(new_n852));
  OAI211_X1 g427(.A(new_n852), .B(KEYINPUT93), .C1(G29), .C2(G32), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n853), .B1(KEYINPUT93), .B2(new_n852), .ZN(new_n854));
  XNOR2_X1  g429(.A(KEYINPUT27), .B(G1996), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(KEYINPUT94), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n854), .B(new_n856), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n826), .A2(new_n828), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT96), .Z(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n769), .A2(new_n770), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n844), .A2(new_n857), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT28), .ZN(new_n863));
  INV_X1    g438(.A(G26), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n863), .B1(new_n864), .B2(G29), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(G29), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n482), .A2(G128), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n484), .A2(G140), .ZN(new_n868));
  NOR2_X1   g443(.A1(G104), .A2(G2105), .ZN(new_n869));
  OAI21_X1  g444(.A(G2104), .B1(new_n462), .B2(G116), .ZN(new_n870));
  OAI211_X1 g445(.A(new_n867), .B(new_n868), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n866), .B1(new_n871), .B2(G29), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n865), .B1(new_n872), .B2(new_n863), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(G2067), .ZN(new_n874));
  OAI21_X1  g449(.A(KEYINPUT102), .B1(new_n862), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n861), .ZN(new_n876));
  NOR4_X1   g451(.A1(new_n876), .A2(new_n771), .A3(new_n843), .A4(new_n859), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  INV_X1    g453(.A(new_n874), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n857), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n875), .A2(new_n880), .ZN(G311));
  NAND3_X1  g456(.A1(new_n877), .A2(new_n879), .A3(new_n857), .ZN(G150));
  AOI22_X1  g457(.A1(new_n520), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n883), .A2(new_n531), .ZN(new_n884));
  INV_X1    g459(.A(G55), .ZN(new_n885));
  INV_X1    g460(.A(G93), .ZN(new_n886));
  OAI22_X1  g461(.A1(new_n505), .A2(new_n885), .B1(new_n513), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g462(.A(G860), .B1(new_n884), .B2(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n888), .B(KEYINPUT37), .Z(new_n889));
  NAND2_X1  g464(.A1(new_n624), .A2(G559), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT39), .ZN(new_n891));
  XNOR2_X1  g466(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n891), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n554), .B1(new_n884), .B2(new_n887), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n884), .A2(new_n887), .ZN(new_n895));
  OAI221_X1 g470(.A(new_n551), .B1(new_n552), .B2(new_n513), .C1(new_n549), .C2(new_n531), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(new_n893), .B(new_n898), .Z(new_n899));
  OAI21_X1  g474(.A(new_n889), .B1(new_n899), .B2(G860), .ZN(G145));
  XNOR2_X1  g475(.A(new_n644), .B(new_n871), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n790), .A2(new_n478), .A3(new_n652), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n652), .B1(new_n790), .B2(new_n478), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n488), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n652), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n791), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(G162), .A3(new_n903), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n823), .B(new_n502), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n906), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n911), .B1(new_n906), .B2(new_n909), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n847), .A2(new_n851), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n482), .A2(G130), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n484), .A2(G142), .ZN(new_n917));
  NOR2_X1   g492(.A1(G106), .A2(G2105), .ZN(new_n918));
  OAI21_X1  g493(.A(G2104), .B1(new_n462), .B2(G118), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n916), .B(new_n917), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n915), .B(new_n920), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n921), .B(new_n728), .ZN(new_n922));
  NOR3_X1   g497(.A1(new_n913), .A2(new_n914), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n922), .ZN(new_n924));
  NOR3_X1   g499(.A1(new_n904), .A2(new_n905), .A3(new_n488), .ZN(new_n925));
  AOI21_X1  g500(.A(G162), .B1(new_n908), .B2(new_n903), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n910), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n924), .B1(new_n927), .B2(new_n912), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n902), .B1(new_n923), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G37), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n922), .B1(new_n913), .B2(new_n914), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(new_n924), .A3(new_n912), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(new_n901), .A3(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT104), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n929), .A2(new_n936), .A3(new_n930), .A4(new_n933), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT40), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n935), .A2(KEYINPUT40), .A3(new_n937), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(G395));
  XNOR2_X1  g517(.A(new_n639), .B(new_n898), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT41), .ZN(new_n944));
  NAND2_X1  g519(.A1(G299), .A2(new_n624), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n631), .A2(new_n632), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n618), .A2(new_n619), .A3(new_n621), .A4(new_n623), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n946), .A2(new_n947), .A3(new_n565), .A4(new_n568), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT105), .B1(new_n945), .B2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT105), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n633), .B2(new_n947), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n944), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  AND2_X1   g527(.A1(new_n945), .A2(new_n948), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT41), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n943), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n956), .A2(KEYINPUT106), .ZN(new_n957));
  INV_X1    g532(.A(new_n956), .ZN(new_n958));
  OAI21_X1  g533(.A(KEYINPUT106), .B1(new_n943), .B2(new_n953), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(KEYINPUT42), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT42), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n957), .B(new_n962), .C1(new_n958), .C2(new_n959), .ZN(new_n963));
  NAND2_X1  g538(.A1(G305), .A2(G166), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n756), .A2(G303), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n612), .B(G288), .ZN(new_n967));
  AND3_X1   g542(.A1(new_n966), .A2(KEYINPUT108), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT108), .B1(new_n966), .B2(new_n967), .ZN(new_n969));
  NOR2_X1   g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n967), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n971), .A2(KEYINPUT107), .A3(new_n964), .A4(new_n965), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n966), .B2(new_n967), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n961), .A2(new_n963), .A3(new_n977), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n977), .B1(new_n961), .B2(new_n963), .ZN(new_n979));
  OAI21_X1  g554(.A(G868), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n980), .B1(G868), .B2(new_n895), .ZN(G295));
  OAI21_X1  g556(.A(new_n980), .B1(G868), .B2(new_n895), .ZN(G331));
  INV_X1    g557(.A(new_n546), .ZN(new_n983));
  AOI21_X1  g558(.A(KEYINPUT72), .B1(new_n538), .B2(G651), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(G286), .B1(new_n985), .B2(new_n545), .ZN(new_n986));
  NOR2_X1   g561(.A1(G301), .A2(G168), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n898), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(G286), .A3(new_n545), .ZN(new_n989));
  NAND2_X1  g564(.A1(G301), .A2(G168), .ZN(new_n990));
  NAND4_X1  g565(.A1(new_n989), .A2(new_n990), .A3(new_n894), .A4(new_n897), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n988), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n952), .A2(new_n954), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n988), .A2(new_n953), .A3(new_n991), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n976), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n993), .A2(new_n970), .A3(new_n975), .A4(new_n994), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n930), .A3(new_n997), .ZN(new_n998));
  OR2_X1    g573(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT43), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n992), .A2(KEYINPUT41), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n953), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n992), .B(KEYINPUT41), .C1(new_n949), .C2(new_n951), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n975), .A4(new_n970), .ZN(new_n1004));
  AND3_X1   g579(.A1(new_n996), .A2(new_n1004), .A3(new_n930), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n999), .B(KEYINPUT44), .C1(new_n1000), .C2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n998), .A2(KEYINPUT43), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n996), .A2(new_n1004), .A3(new_n1000), .A4(new_n930), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT109), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT109), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n1012), .B(KEYINPUT44), .C1(new_n1007), .C2(new_n1008), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1006), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(KEYINPUT110), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT110), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1016), .B(new_n1006), .C1(new_n1011), .C2(new_n1013), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(G397));
  NOR2_X1   g593(.A1(new_n871), .A2(G2067), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n915), .B(G1996), .ZN(new_n1020));
  XOR2_X1   g595(.A(new_n871), .B(G2067), .Z(new_n1021));
  INV_X1    g596(.A(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n728), .A2(new_n730), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n1019), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(G1384), .B1(new_n494), .B2(new_n501), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(KEYINPUT111), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(KEYINPUT111), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n477), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n471), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n1033));
  OAI211_X1 g608(.A(G40), .B(new_n1032), .C1(new_n1033), .C2(new_n462), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1031), .A2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1025), .A2(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(G290), .A2(G1986), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1040), .B(KEYINPUT48), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1036), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n728), .A2(new_n730), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1024), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1023), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1041), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1036), .A2(G1996), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT46), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(KEYINPUT126), .ZN(new_n1049));
  XNOR2_X1  g624(.A(new_n1047), .B(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(KEYINPUT126), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1022), .A2(new_n915), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1051), .B1(new_n1036), .B2(new_n1052), .ZN(new_n1053));
  OR3_X1    g628(.A1(new_n1050), .A2(KEYINPUT47), .A3(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(KEYINPUT47), .B1(new_n1050), .B2(new_n1053), .ZN(new_n1055));
  AOI211_X1 g630(.A(new_n1037), .B(new_n1046), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(G1384), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n502), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1058), .A2(new_n1034), .ZN(new_n1059));
  INV_X1    g634(.A(G8), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1976), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1062), .B2(G288), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT52), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1063), .A2(KEYINPUT113), .A3(KEYINPUT52), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1063), .A2(KEYINPUT52), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(G1976), .B2(new_n742), .ZN(new_n1070));
  OR3_X1    g645(.A1(G305), .A2(KEYINPUT114), .A3(G1981), .ZN(new_n1071));
  OAI21_X1  g646(.A(KEYINPUT114), .B1(G305), .B2(G1981), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(new_n598), .B(KEYINPUT115), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1074), .A2(new_n753), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G1981), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1073), .A2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT49), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1077), .A2(KEYINPUT116), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT116), .ZN(new_n1080));
  OAI211_X1 g655(.A(new_n1073), .B(new_n1076), .C1(new_n1080), .C2(KEYINPUT49), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1079), .A2(new_n1061), .A3(new_n1081), .ZN(new_n1082));
  AND3_X1   g657(.A1(new_n1068), .A2(new_n1070), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1034), .B1(new_n1058), .B2(new_n1028), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1026), .A2(KEYINPUT45), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1971), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT50), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1058), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1026), .A2(KEYINPUT50), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1034), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(G2090), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1060), .B1(new_n1088), .B2(new_n1094), .ZN(new_n1095));
  NOR2_X1   g670(.A1(G166), .A2(new_n1060), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT55), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT112), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT112), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1095), .A2(new_n1100), .A3(new_n1097), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1085), .A2(KEYINPUT118), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1026), .A2(new_n1104), .A3(KEYINPUT45), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1084), .A2(new_n1103), .A3(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n828), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1092), .A2(new_n793), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1060), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1109), .A2(G168), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1110), .A2(new_n1111), .A3(KEYINPUT63), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1083), .B1(new_n1102), .B2(new_n1112), .ZN(new_n1113));
  OR2_X1    g688(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1068), .A2(new_n1070), .A3(new_n1082), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT63), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  XOR2_X1   g691(.A(new_n1061), .B(KEYINPUT117), .Z(new_n1117));
  AND3_X1   g692(.A1(new_n1082), .A2(new_n1062), .A3(new_n742), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1073), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1117), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1113), .A2(new_n1116), .A3(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(G168), .A2(new_n1060), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT51), .B1(new_n1123), .B2(KEYINPUT123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1124), .B1(new_n1109), .B2(new_n1122), .ZN(new_n1125));
  AOI22_X1  g700(.A1(new_n1106), .A2(new_n828), .B1(new_n1092), .B2(new_n793), .ZN(new_n1126));
  OAI221_X1 g701(.A(new_n1123), .B1(KEYINPUT123), .B2(KEYINPUT51), .C1(new_n1126), .C2(new_n1060), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1109), .A2(G286), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1058), .A2(new_n1028), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1130), .A2(new_n817), .A3(new_n1085), .A4(new_n1035), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT53), .ZN(new_n1132));
  AOI21_X1  g707(.A(KEYINPUT50), .B1(new_n502), .B2(new_n1057), .ZN(new_n1133));
  AOI211_X1 g708(.A(new_n1089), .B(G1384), .C1(new_n494), .C2(new_n501), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1035), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1131), .A2(new_n1132), .B1(new_n1135), .B2(new_n788), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n1132), .A2(G2078), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1084), .A2(new_n1103), .A3(new_n1105), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(G171), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1129), .B1(KEYINPUT62), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1135), .A2(new_n774), .ZN(new_n1143));
  NOR3_X1   g718(.A1(new_n1058), .A2(new_n1034), .A3(G2067), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n947), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(G1956), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1135), .A2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT119), .B(G2072), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT56), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1130), .A2(new_n1085), .A3(new_n1035), .A4(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n633), .B(KEYINPUT57), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1148), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1146), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1152), .B1(new_n1148), .B2(new_n1151), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1155), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1154), .A2(KEYINPUT120), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT120), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  XOR2_X1   g734(.A(KEYINPUT121), .B(G1996), .Z(new_n1160));
  NAND4_X1  g735(.A1(new_n1130), .A2(new_n1085), .A3(new_n1035), .A4(new_n1160), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT58), .B(G1341), .Z(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(new_n1058), .B2(new_n1034), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  AOI22_X1  g739(.A1(new_n1164), .A2(new_n554), .B1(KEYINPUT122), .B2(KEYINPUT59), .ZN(new_n1165));
  NAND2_X1  g740(.A1(KEYINPUT122), .A2(KEYINPUT59), .ZN(new_n1166));
  AOI211_X1 g741(.A(new_n896), .B(new_n1166), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n947), .A2(KEYINPUT60), .ZN(new_n1168));
  AOI211_X1 g743(.A(new_n1168), .B(new_n1144), .C1(new_n774), .C2(new_n1135), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1165), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1170));
  AOI211_X1 g745(.A(new_n624), .B(new_n1144), .C1(new_n774), .C2(new_n1135), .ZN(new_n1171));
  OAI21_X1  g746(.A(KEYINPUT60), .B1(new_n1171), .B2(new_n1146), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT61), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1153), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1173), .B1(new_n1174), .B2(new_n1155), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1156), .A2(KEYINPUT61), .A3(new_n1153), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1170), .A2(new_n1172), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1159), .A2(new_n1177), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1030), .A2(new_n1085), .A3(new_n1035), .A4(new_n1137), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1136), .A2(new_n1179), .A3(G301), .ZN(new_n1180));
  AOI21_X1  g755(.A(KEYINPUT54), .B1(new_n1140), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT125), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1136), .A2(new_n1179), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1182), .B1(new_n1183), .B2(G171), .ZN(new_n1184));
  AOI211_X1 g759(.A(KEYINPUT125), .B(G301), .C1(new_n1136), .C2(new_n1179), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(KEYINPUT54), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1139), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1187), .B1(new_n1188), .B2(G301), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1181), .B1(new_n1186), .B2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1178), .A2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1129), .A2(KEYINPUT62), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1192), .A2(new_n1141), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1142), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1111), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1195));
  AND3_X1   g770(.A1(new_n1083), .A2(new_n1195), .A3(KEYINPUT124), .ZN(new_n1196));
  AOI21_X1  g771(.A(KEYINPUT124), .B1(new_n1083), .B2(new_n1195), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1121), .B1(new_n1194), .B2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1045), .B1(G1986), .B2(G290), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1036), .B1(new_n1200), .B2(new_n1039), .ZN(new_n1201));
  OAI21_X1  g776(.A(new_n1056), .B1(new_n1199), .B2(new_n1201), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g777(.A(G227), .ZN(new_n1204));
  AND2_X1   g778(.A1(new_n674), .A2(new_n460), .ZN(new_n1205));
  NAND4_X1  g779(.A1(new_n719), .A2(new_n722), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n1206), .A2(KEYINPUT127), .ZN(new_n1207));
  NAND2_X1  g781(.A1(new_n1207), .A2(new_n1009), .ZN(new_n1208));
  OAI21_X1  g782(.A(new_n934), .B1(new_n1206), .B2(KEYINPUT127), .ZN(new_n1209));
  NOR2_X1   g783(.A1(new_n1208), .A2(new_n1209), .ZN(G308));
  OR2_X1    g784(.A1(new_n1206), .A2(KEYINPUT127), .ZN(new_n1211));
  NAND4_X1  g785(.A1(new_n1211), .A2(new_n934), .A3(new_n1009), .A4(new_n1207), .ZN(G225));
endmodule


