//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 0 0 1 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n243, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1270, new_n1272, new_n1273,
    new_n1274, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1344, new_n1345;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n210), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  OR2_X1    g0019(.A1(new_n219), .A2(KEYINPUT0), .ZN(new_n220));
  OAI21_X1  g0020(.A(G50), .B1(G58), .B2(G68), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(G20), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n219), .A2(KEYINPUT0), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n220), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT66), .Z(new_n228));
  INV_X1    g0028(.A(G68), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(KEYINPUT67), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT67), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n231), .A2(G68), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(G238), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI22_X1  g0036(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n237));
  AOI22_X1  g0037(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n238));
  AOI22_X1  g0038(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n239));
  NAND2_X1  g0039(.A1(G58), .A2(G232), .ZN(new_n240));
  NAND4_X1  g0040(.A1(new_n237), .A2(new_n238), .A3(new_n239), .A4(new_n240), .ZN(new_n241));
  OAI21_X1  g0041(.A(new_n214), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT1), .ZN(new_n243));
  NOR2_X1   g0043(.A1(new_n228), .A2(new_n243), .ZN(G361));
  XOR2_X1   g0044(.A(G238), .B(G244), .Z(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT68), .B(KEYINPUT2), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G226), .B(G232), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G250), .B(G257), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G264), .B(G270), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G358));
  XNOR2_X1  g0053(.A(G87), .B(G97), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G107), .B(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(G50), .B(G68), .ZN(new_n257));
  XNOR2_X1  g0057(.A(G58), .B(G77), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n256), .B(new_n259), .ZN(G351));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n223), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(KEYINPUT70), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT70), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n264), .B1(new_n261), .B2(new_n223), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G13), .ZN(new_n268));
  NOR3_X1   g0068(.A1(new_n268), .A2(new_n212), .A3(G1), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n211), .A2(G20), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n270), .A2(G50), .A3(new_n271), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n212), .B1(new_n201), .B2(new_n202), .ZN(new_n273));
  NOR2_X1   g0073(.A1(G20), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G150), .ZN(new_n275));
  XNOR2_X1  g0075(.A(KEYINPUT8), .B(G58), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n212), .A2(G33), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n267), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n269), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n272), .B(new_n279), .C1(G50), .C2(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(new_n281), .B(KEYINPUT9), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT69), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G41), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n211), .B(G274), .C1(new_n287), .C2(G45), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n223), .B1(G33), .B2(G41), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n289), .B1(G226), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT3), .B(G33), .ZN(new_n296));
  NOR2_X1   g0096(.A1(G222), .A2(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(G1698), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(G223), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n296), .B1(new_n297), .B2(new_n299), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n300), .B(new_n290), .C1(G77), .C2(new_n296), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G190), .ZN(new_n304));
  INV_X1    g0104(.A(G200), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n282), .B(new_n304), .C1(new_n305), .C2(new_n303), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT10), .ZN(new_n307));
  INV_X1    g0107(.A(G179), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n302), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n281), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(G33), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(KEYINPUT3), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT3), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(G33), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n317), .A3(KEYINPUT74), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT74), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n319), .A2(new_n314), .A3(KEYINPUT3), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  MUX2_X1   g0121(.A(G223), .B(G226), .S(G1698), .Z(new_n322));
  AOI22_X1  g0122(.A1(new_n321), .A2(new_n322), .B1(G33), .B2(G87), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n323), .A2(new_n291), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n289), .B1(G232), .B2(new_n294), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(new_n308), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(G169), .B2(new_n326), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G58), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n230), .B2(new_n232), .ZN(new_n331));
  OAI21_X1  g0131(.A(G20), .B1(new_n331), .B2(new_n201), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT76), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n274), .A2(G159), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n333), .B1(new_n332), .B2(new_n334), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT78), .B1(new_n316), .B2(G33), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT78), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n339), .A2(new_n314), .A3(KEYINPUT3), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n338), .A2(new_n340), .A3(new_n317), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT7), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n342), .A2(G20), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n342), .B1(new_n296), .B2(G20), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n234), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n336), .A2(new_n337), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n262), .B1(new_n347), .B2(KEYINPUT16), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n321), .A2(KEYINPUT75), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT75), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n318), .A2(new_n320), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n349), .A2(new_n212), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n342), .ZN(new_n353));
  NOR3_X1   g0153(.A1(new_n316), .A2(KEYINPUT74), .A3(G33), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n296), .B2(KEYINPUT74), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n343), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n229), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n337), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n358), .A2(new_n335), .A3(KEYINPUT16), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT77), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT16), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n336), .A2(new_n337), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT77), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n352), .A2(new_n342), .B1(new_n355), .B2(new_n343), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n362), .B(new_n363), .C1(new_n229), .C2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n348), .B1(new_n360), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(new_n276), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n270), .A2(new_n367), .A3(new_n271), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n280), .B2(new_n367), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n329), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT18), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT18), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(new_n329), .C1(new_n366), .C2(new_n369), .ZN(new_n373));
  XNOR2_X1  g0173(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n360), .A2(new_n365), .ZN(new_n375));
  INV_X1    g0175(.A(new_n348), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n369), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n326), .A2(G190), .ZN(new_n378));
  AOI21_X1  g0178(.A(G200), .B1(new_n324), .B2(new_n325), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n374), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT17), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(KEYINPUT79), .ZN(new_n384));
  NOR4_X1   g0184(.A1(new_n366), .A2(new_n369), .A3(new_n380), .A4(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n371), .B(new_n373), .C1(new_n382), .C2(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n288), .B1(new_n293), .B2(new_n235), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n298), .A2(G232), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n296), .B(new_n388), .C1(G226), .C2(G1698), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G97), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n291), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  XNOR2_X1  g0192(.A(KEYINPUT72), .B(KEYINPUT13), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n394), .A2(G169), .ZN(new_n395));
  MUX2_X1   g0195(.A(KEYINPUT13), .B(new_n393), .S(new_n392), .Z(new_n396));
  OAI22_X1  g0196(.A1(new_n395), .A2(KEYINPUT14), .B1(new_n396), .B2(new_n308), .ZN(new_n397));
  AND2_X1   g0197(.A1(new_n395), .A2(KEYINPUT14), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n274), .A2(G50), .ZN(new_n399));
  OAI221_X1 g0199(.A(new_n399), .B1(new_n203), .B2(new_n277), .C1(new_n233), .C2(new_n212), .ZN(new_n400));
  AOI21_X1  g0200(.A(KEYINPUT11), .B1(new_n267), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n267), .A2(KEYINPUT11), .A3(new_n400), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n269), .A2(new_n262), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(G68), .A3(new_n271), .ZN(new_n404));
  OR3_X1    g0204(.A1(new_n280), .A2(KEYINPUT12), .A3(G68), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT73), .ZN(new_n406));
  OAI21_X1  g0206(.A(KEYINPUT12), .B1(new_n280), .B2(new_n233), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g0208(.A1(new_n405), .A2(KEYINPUT73), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n402), .B(new_n404), .C1(new_n408), .C2(new_n409), .ZN(new_n410));
  OAI22_X1  g0210(.A1(new_n397), .A2(new_n398), .B1(new_n401), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n394), .A2(G200), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n410), .A2(new_n401), .ZN(new_n413));
  INV_X1    g0213(.A(G190), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n412), .B(new_n413), .C1(new_n396), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n411), .A2(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  XOR2_X1   g0217(.A(new_n276), .B(KEYINPUT71), .Z(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n274), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT15), .B(G87), .ZN(new_n420));
  OAI221_X1 g0220(.A(new_n419), .B1(new_n212), .B2(new_n203), .C1(new_n277), .C2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n262), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n203), .B1(new_n211), .B2(G20), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n403), .A2(new_n423), .B1(new_n203), .B2(new_n269), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n296), .A2(G232), .A3(new_n298), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(new_n207), .B2(new_n296), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n315), .A2(new_n317), .ZN(new_n428));
  NOR3_X1   g0228(.A1(new_n428), .A2(new_n235), .A3(new_n298), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n290), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(G244), .ZN(new_n431));
  OAI211_X1 g0231(.A(new_n430), .B(new_n288), .C1(new_n431), .C2(new_n293), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(G200), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n425), .B(new_n433), .C1(new_n414), .C2(new_n432), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n422), .A2(new_n424), .B1(new_n310), .B2(new_n432), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n432), .A2(G179), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g0237(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n417), .A2(new_n438), .ZN(new_n439));
  NOR3_X1   g0239(.A1(new_n313), .A2(new_n386), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT81), .ZN(new_n442));
  INV_X1    g0242(.A(G45), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G1), .ZN(new_n444));
  XNOR2_X1  g0244(.A(KEYINPUT69), .B(G41), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n442), .B(new_n444), .C1(new_n445), .C2(KEYINPUT5), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n283), .A2(KEYINPUT5), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT5), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n285), .A2(G41), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n283), .A2(KEYINPUT69), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n449), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n442), .B1(new_n452), .B2(new_n444), .ZN(new_n453));
  OAI211_X1 g0253(.A(G264), .B(new_n291), .C1(new_n448), .C2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT90), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT5), .B1(new_n284), .B2(new_n286), .ZN(new_n456));
  INV_X1    g0256(.A(new_n444), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT81), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n458), .A2(new_n447), .A3(new_n446), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT90), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(G264), .A4(new_n291), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n455), .A2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(G274), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n290), .A2(new_n463), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n458), .A2(new_n447), .A3(new_n446), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n217), .A2(G1698), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n321), .B(new_n466), .C1(G250), .C2(G1698), .ZN(new_n467));
  INV_X1    g0267(.A(G294), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n314), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n291), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n462), .A2(new_n414), .A3(new_n465), .A4(new_n472), .ZN(new_n473));
  AND4_X1   g0273(.A1(new_n458), .A2(new_n447), .A3(new_n446), .A4(new_n464), .ZN(new_n474));
  AOI211_X1 g0274(.A(new_n474), .B(new_n471), .C1(new_n455), .C2(new_n461), .ZN(new_n475));
  OAI211_X1 g0275(.A(new_n473), .B(KEYINPUT91), .C1(new_n475), .C2(G200), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n462), .A2(new_n465), .A3(new_n472), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT91), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(new_n305), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT24), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT87), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT22), .ZN(new_n482));
  AOI21_X1  g0282(.A(G20), .B1(new_n318), .B2(new_n320), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n482), .B1(new_n483), .B2(G87), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n482), .A2(new_n212), .A3(G87), .ZN(new_n485));
  OAI21_X1  g0285(.A(KEYINPUT86), .B1(new_n428), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT86), .ZN(new_n487));
  INV_X1    g0287(.A(G87), .ZN(new_n488));
  NOR3_X1   g0288(.A1(new_n488), .A2(KEYINPUT22), .A3(G20), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n296), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n481), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n428), .A2(KEYINPUT86), .A3(new_n485), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n487), .B1(new_n296), .B2(new_n489), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI211_X1 g0295(.A(G20), .B(new_n488), .C1(new_n318), .C2(new_n320), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n495), .B(KEYINPUT87), .C1(new_n496), .C2(new_n482), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  OR3_X1    g0298(.A1(new_n212), .A2(KEYINPUT23), .A3(G107), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n212), .A2(G33), .A3(G116), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT88), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT23), .B1(new_n212), .B2(G107), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n499), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n502), .A2(new_n501), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n480), .B1(new_n498), .B2(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n505), .ZN(new_n507));
  AOI211_X1 g0307(.A(KEYINPUT24), .B(new_n507), .C1(new_n492), .C2(new_n497), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n262), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT25), .ZN(new_n510));
  AOI211_X1 g0310(.A(G107), .B(new_n280), .C1(KEYINPUT89), .C2(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n510), .A2(KEYINPUT89), .ZN(new_n512));
  XOR2_X1   g0312(.A(new_n511), .B(new_n512), .Z(new_n513));
  NOR2_X1   g0313(.A1(new_n314), .A2(G1), .ZN(new_n514));
  NOR4_X1   g0314(.A1(new_n263), .A2(new_n265), .A3(new_n269), .A4(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n516), .A2(new_n207), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  NAND4_X1  g0318(.A1(new_n476), .A2(new_n479), .A3(new_n509), .A4(new_n518), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n462), .A2(new_n308), .A3(new_n465), .A4(new_n472), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n475), .B2(G169), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n509), .A2(new_n518), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n519), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n207), .B1(new_n344), .B2(new_n345), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n274), .A2(G77), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n207), .A2(KEYINPUT6), .A3(G97), .ZN(new_n528));
  XNOR2_X1  g0328(.A(G97), .B(G107), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT6), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n527), .B1(new_n531), .B2(new_n212), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n262), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n280), .A2(G97), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n534), .B1(new_n515), .B2(G97), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT80), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n533), .A2(KEYINPUT80), .A3(new_n535), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n431), .B1(new_n318), .B2(new_n320), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT4), .B1(new_n541), .B2(new_n298), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n315), .A2(new_n317), .A3(G250), .A4(G1698), .ZN(new_n543));
  AND2_X1   g0343(.A1(KEYINPUT4), .A2(G244), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n315), .A2(new_n317), .A3(new_n544), .A4(new_n298), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G283), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n290), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n459), .A2(G257), .A3(new_n291), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n548), .A2(new_n549), .A3(new_n414), .A4(new_n465), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(new_n465), .A3(new_n549), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n305), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n540), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n515), .A2(G87), .ZN(new_n554));
  INV_X1    g0354(.A(new_n262), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n321), .A2(new_n212), .A3(G68), .ZN(new_n556));
  NOR3_X1   g0356(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n557));
  AOI21_X1  g0357(.A(G20), .B1(G33), .B2(G97), .ZN(new_n558));
  OAI21_X1  g0358(.A(KEYINPUT19), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n560), .A2(new_n212), .A3(G33), .A4(G97), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n555), .B1(new_n556), .B2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT82), .ZN(new_n564));
  INV_X1    g0364(.A(new_n420), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n280), .ZN(new_n566));
  NOR3_X1   g0366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  AOI211_X1 g0367(.A(G20), .B(new_n229), .C1(new_n318), .C2(new_n320), .ZN(new_n568));
  AND2_X1   g0368(.A1(new_n559), .A2(new_n561), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n262), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n566), .ZN(new_n571));
  AOI21_X1  g0371(.A(KEYINPUT82), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n554), .B1(new_n567), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n235), .A2(G1698), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n321), .A2(new_n574), .B1(G33), .B2(G116), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n541), .A2(G1698), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n291), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n457), .A2(new_n210), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n444), .A2(new_n463), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n578), .A2(new_n291), .A3(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g0381(.A(G200), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n574), .ZN(new_n583));
  INV_X1    g0383(.A(G116), .ZN(new_n584));
  OAI22_X1  g0384(.A1(new_n355), .A2(new_n583), .B1(new_n314), .B2(new_n584), .ZN(new_n585));
  AOI211_X1 g0385(.A(new_n431), .B(new_n298), .C1(new_n318), .C2(new_n320), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n290), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n587), .A2(G190), .A3(new_n580), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n564), .B1(new_n563), .B2(new_n566), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n570), .A2(KEYINPUT82), .A3(new_n571), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n590), .A2(new_n591), .B1(new_n515), .B2(new_n565), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n310), .B1(new_n577), .B2(new_n581), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n587), .A2(new_n308), .A3(new_n580), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  OAI22_X1  g0395(.A1(new_n573), .A2(new_n589), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n551), .A2(G169), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n548), .A2(new_n549), .A3(G179), .A4(new_n465), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n597), .A2(new_n598), .B1(new_n533), .B2(new_n535), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n553), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n459), .A2(G270), .A3(new_n291), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n218), .A2(G1698), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(G257), .B2(G1698), .ZN(new_n603));
  INV_X1    g0403(.A(G303), .ZN(new_n604));
  OAI22_X1  g0404(.A1(new_n355), .A2(new_n603), .B1(new_n604), .B2(new_n296), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n290), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n601), .A2(new_n465), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(G200), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n514), .A2(new_n584), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n268), .A2(G1), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n212), .A2(G116), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n403), .A2(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI211_X1 g0412(.A(new_n546), .B(new_n212), .C1(G33), .C2(new_n206), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n613), .B(new_n262), .C1(new_n212), .C2(G116), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT20), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n612), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n608), .B(new_n619), .C1(new_n414), .C2(new_n607), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT85), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n618), .A2(G169), .ZN(new_n622));
  AOI21_X1  g0422(.A(KEYINPUT21), .B1(new_n622), .B2(new_n607), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n308), .B1(new_n605), .B2(new_n290), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(new_n601), .A3(new_n465), .ZN(new_n625));
  OAI21_X1  g0425(.A(KEYINPUT84), .B1(new_n625), .B2(new_n619), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n601), .A2(new_n624), .A3(new_n465), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT84), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n628), .A3(new_n618), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n623), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n607), .A2(KEYINPUT21), .A3(G169), .A4(new_n618), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT83), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n622), .A2(KEYINPUT83), .A3(KEYINPUT21), .A4(new_n607), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n600), .A2(new_n621), .A3(new_n636), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n441), .A2(new_n525), .A3(new_n637), .ZN(G372));
  INV_X1    g0438(.A(new_n312), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n411), .A2(new_n437), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n640), .B(new_n415), .C1(new_n382), .C2(new_n385), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n371), .A2(new_n373), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n639), .B1(new_n643), .B2(new_n307), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  INV_X1    g0445(.A(new_n595), .ZN(new_n646));
  OAI22_X1  g0446(.A1(new_n567), .A2(new_n572), .B1(new_n516), .B2(new_n420), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n590), .A2(new_n591), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n649), .A2(new_n554), .A3(new_n582), .A4(new_n588), .ZN(new_n650));
  AOI22_X1  g0450(.A1(new_n597), .A2(new_n598), .B1(new_n538), .B2(new_n539), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n648), .B(new_n650), .C1(new_n651), .C2(KEYINPUT92), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n597), .A2(new_n598), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n653), .A2(KEYINPUT92), .A3(new_n540), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n645), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n596), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(KEYINPUT26), .A3(new_n599), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n521), .B1(new_n509), .B2(new_n518), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n630), .A2(new_n635), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n600), .B(new_n519), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n658), .A2(new_n661), .A3(new_n648), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n644), .B1(new_n441), .B2(new_n663), .ZN(G369));
  AND2_X1   g0464(.A1(new_n621), .A2(new_n636), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n610), .A2(new_n212), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(KEYINPUT27), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(G213), .A3(new_n668), .ZN(new_n669));
  XOR2_X1   g0469(.A(KEYINPUT93), .B(G343), .Z(new_n670));
  NOR2_X1   g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n619), .A2(new_n672), .ZN(new_n673));
  MUX2_X1   g0473(.A(new_n665), .B(new_n660), .S(new_n673), .Z(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n513), .A2(new_n517), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n507), .B1(new_n492), .B2(new_n497), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n678), .B(new_n480), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n677), .B1(new_n679), .B2(new_n262), .ZN(new_n680));
  OAI21_X1  g0480(.A(KEYINPUT94), .B1(new_n680), .B2(new_n672), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT94), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n523), .A2(new_n682), .A3(new_n671), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n681), .A2(new_n519), .A3(new_n524), .A4(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT95), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n519), .A2(new_n524), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n687), .A2(KEYINPUT95), .A3(new_n683), .A4(new_n681), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n524), .A2(new_n672), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n676), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n636), .A2(new_n671), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n686), .A2(new_n688), .A3(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT96), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n659), .A2(new_n672), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n696), .B1(new_n695), .B2(new_n697), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n693), .B1(new_n698), .B2(new_n699), .ZN(G399));
  NOR2_X1   g0500(.A1(new_n216), .A2(new_n287), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NOR3_X1   g0502(.A1(new_n208), .A2(G87), .A3(G116), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n702), .A2(G1), .A3(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n222), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n705), .B2(new_n702), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n663), .A2(KEYINPUT29), .A3(new_n671), .ZN(new_n708));
  INV_X1    g0508(.A(new_n648), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n552), .A2(new_n550), .ZN(new_n710));
  INV_X1    g0510(.A(new_n539), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT80), .B1(new_n533), .B2(new_n535), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n547), .ZN(new_n715));
  AOI211_X1 g0515(.A(new_n431), .B(G1698), .C1(new_n318), .C2(new_n320), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(KEYINPUT4), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n474), .B1(new_n290), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n310), .B1(new_n718), .B2(new_n549), .ZN(new_n719));
  INV_X1    g0519(.A(new_n598), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n536), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n714), .A2(new_n721), .A3(new_n648), .A4(new_n650), .ZN(new_n722));
  AND3_X1   g0522(.A1(new_n479), .A2(new_n509), .A3(new_n518), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n476), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n636), .A2(new_n524), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n709), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n596), .A2(new_n721), .A3(KEYINPUT26), .ZN(new_n727));
  INV_X1    g0527(.A(new_n654), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n651), .A2(KEYINPUT92), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n728), .A2(new_n729), .A3(new_n656), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n727), .B1(new_n730), .B2(KEYINPUT26), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n671), .B1(new_n726), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(G330), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n665), .A2(new_n687), .A3(new_n600), .A4(new_n672), .ZN(new_n736));
  AOI21_X1  g0536(.A(G179), .B1(new_n587), .B2(new_n580), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT97), .ZN(new_n738));
  AND3_X1   g0538(.A1(new_n737), .A2(new_n738), .A3(new_n607), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n738), .B1(new_n737), .B2(new_n607), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n477), .B(new_n551), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n587), .A2(new_n580), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n551), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n471), .B1(new_n455), .B2(new_n461), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n743), .A2(new_n744), .A3(new_n627), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT30), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n743), .A2(KEYINPUT30), .A3(new_n744), .A4(new_n627), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n741), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n671), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  AOI21_X1  g0551(.A(KEYINPUT31), .B1(new_n749), .B2(new_n671), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n735), .B1(new_n736), .B2(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n708), .A2(new_n734), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n707), .B1(new_n755), .B2(G1), .ZN(G364));
  NOR2_X1   g0556(.A1(new_n268), .A2(G20), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n211), .B1(new_n757), .B2(G45), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n702), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n676), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n761), .B1(G330), .B2(new_n674), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n215), .A2(new_n296), .ZN(new_n763));
  INV_X1    g0563(.A(G355), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n763), .A2(new_n764), .B1(G116), .B2(new_n215), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n705), .A2(G45), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(G45), .B2(new_n259), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n349), .A2(new_n351), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n216), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n765), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n223), .B1(G20), .B2(new_n310), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n760), .B1(new_n770), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n212), .A2(new_n308), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G190), .A2(G200), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(G311), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n212), .A2(G179), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n779), .ZN(new_n783));
  INV_X1    g0583(.A(G329), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n780), .A2(new_n781), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n778), .A2(G190), .A3(new_n305), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n296), .B(new_n785), .C1(G322), .C2(new_n787), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n782), .A2(new_n414), .A3(G200), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT98), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G283), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n778), .A2(G200), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n414), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n782), .A2(G190), .A3(G200), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n793), .A2(G326), .B1(new_n795), .B2(G303), .ZN(new_n796));
  NOR3_X1   g0596(.A1(new_n414), .A2(G179), .A3(G200), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n797), .A2(new_n212), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n792), .A2(G190), .ZN(new_n800));
  XNOR2_X1  g0600(.A(KEYINPUT33), .B(G317), .ZN(new_n801));
  AOI22_X1  g0601(.A1(G294), .A2(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n788), .A2(new_n791), .A3(new_n796), .A4(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT99), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n800), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n806), .A2(new_n229), .B1(new_n794), .B2(new_n488), .ZN(new_n807));
  INV_X1    g0607(.A(new_n793), .ZN(new_n808));
  INV_X1    g0608(.A(new_n783), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(G159), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n808), .A2(new_n202), .B1(new_n810), .B2(KEYINPUT32), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n807), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n790), .A2(G107), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n296), .B1(new_n786), .B2(new_n330), .ZN(new_n814));
  INV_X1    g0614(.A(new_n780), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(G77), .B2(new_n815), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n810), .A2(KEYINPUT32), .B1(new_n799), .B2(G97), .ZN(new_n817));
  NAND4_X1  g0617(.A1(new_n812), .A2(new_n813), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n803), .A2(new_n804), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n805), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n777), .B1(new_n820), .B2(new_n774), .ZN(new_n821));
  INV_X1    g0621(.A(new_n773), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n674), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n762), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(G396));
  INV_X1    g0625(.A(new_n774), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n772), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n799), .A2(G97), .B1(new_n795), .B2(G107), .ZN(new_n828));
  INV_X1    g0628(.A(G283), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n829), .B2(new_n806), .C1(new_n604), .C2(new_n808), .ZN(new_n830));
  INV_X1    g0630(.A(new_n790), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(new_n488), .ZN(new_n832));
  AOI22_X1  g0632(.A1(new_n787), .A2(G294), .B1(new_n809), .B2(G311), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n833), .B(new_n428), .C1(new_n584), .C2(new_n780), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n830), .A2(new_n832), .A3(new_n834), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n787), .A2(G143), .B1(new_n815), .B2(G159), .ZN(new_n836));
  INV_X1    g0636(.A(G137), .ZN(new_n837));
  INV_X1    g0637(.A(G150), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n836), .B1(new_n808), .B2(new_n837), .C1(new_n838), .C2(new_n806), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT34), .ZN(new_n840));
  INV_X1    g0640(.A(new_n768), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n799), .A2(G58), .B1(G132), .B2(new_n809), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n202), .B2(new_n794), .ZN(new_n843));
  AOI211_X1 g0643(.A(new_n841), .B(new_n843), .C1(G68), .C2(new_n790), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n835), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n760), .B1(G77), .B2(new_n827), .C1(new_n845), .C2(new_n826), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n434), .B1(new_n425), .B2(new_n672), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(new_n437), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n435), .A2(new_n436), .A3(new_n672), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n846), .B1(new_n850), .B2(new_n771), .ZN(new_n851));
  XOR2_X1   g0651(.A(new_n851), .B(KEYINPUT100), .Z(new_n852));
  AND2_X1   g0652(.A1(new_n438), .A2(new_n672), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n662), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT101), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n662), .A2(KEYINPUT101), .A3(new_n853), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n850), .B1(new_n663), .B2(new_n671), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n754), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(new_n760), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n858), .A2(new_n754), .A3(new_n859), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n852), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(G384));
  NOR2_X1   g0664(.A1(new_n757), .A2(new_n211), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT40), .ZN(new_n866));
  INV_X1    g0666(.A(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n375), .A2(new_n376), .ZN(new_n868));
  INV_X1    g0668(.A(new_n369), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n868), .A2(new_n869), .A3(new_n381), .ZN(new_n870));
  INV_X1    g0670(.A(new_n669), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n871), .B1(new_n366), .B2(new_n369), .ZN(new_n872));
  XNOR2_X1  g0672(.A(KEYINPUT104), .B(KEYINPUT37), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n870), .A2(new_n370), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  OAI211_X1 g0674(.A(new_n335), .B(new_n358), .C1(new_n364), .C2(new_n229), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n266), .B1(new_n875), .B2(new_n361), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n375), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n328), .B1(new_n877), .B2(new_n869), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n669), .B1(new_n877), .B2(new_n869), .ZN(new_n879));
  NOR3_X1   g0679(.A1(new_n366), .A2(new_n369), .A3(new_n380), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT37), .ZN(new_n882));
  OAI211_X1 g0682(.A(KEYINPUT105), .B(new_n874), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n386), .A2(new_n879), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n877), .A2(new_n869), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n871), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n870), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT37), .B1(new_n888), .B2(new_n878), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT105), .B1(new_n889), .B2(new_n874), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n867), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT105), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n886), .A2(new_n871), .B1(new_n377), .B2(new_n381), .ZN(new_n893));
  INV_X1    g0693(.A(new_n878), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n882), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n874), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n892), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n897), .A2(KEYINPUT38), .A3(new_n883), .A4(new_n884), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n891), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT107), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n637), .A2(new_n525), .A3(new_n671), .ZN(new_n901));
  INV_X1    g0701(.A(new_n752), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n750), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n900), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n413), .A2(new_n672), .ZN(new_n905));
  OR2_X1    g0705(.A1(new_n416), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n416), .A2(new_n905), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n850), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n736), .A2(new_n753), .A3(KEYINPUT107), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n904), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n866), .B1(new_n899), .B2(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(new_n872), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n386), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n870), .A2(new_n370), .A3(new_n872), .ZN(new_n914));
  INV_X1    g0714(.A(new_n873), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g0716(.A1(new_n916), .A2(new_n874), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n867), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n898), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT108), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n898), .A2(new_n918), .A3(KEYINPUT108), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n904), .A2(new_n908), .A3(new_n909), .A4(KEYINPUT40), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n921), .A2(new_n922), .A3(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n911), .A2(new_n925), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n440), .A2(new_n904), .A3(new_n909), .ZN(new_n927));
  OAI21_X1  g0727(.A(G330), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n928), .A2(KEYINPUT109), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(KEYINPUT109), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n926), .A2(new_n927), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT39), .B1(new_n898), .B2(new_n918), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n891), .A2(KEYINPUT39), .A3(new_n898), .ZN(new_n935));
  OR3_X1    g0735(.A1(new_n411), .A2(KEYINPUT106), .A3(new_n671), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT106), .B1(new_n411), .B2(new_n671), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n934), .A2(new_n935), .A3(new_n938), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n642), .A2(new_n871), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT103), .ZN(new_n942));
  AND3_X1   g0742(.A1(new_n662), .A2(KEYINPUT101), .A3(new_n853), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT101), .B1(new_n662), .B2(new_n853), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n849), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n906), .A2(new_n907), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n899), .B1(new_n942), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n945), .A2(KEYINPUT103), .A3(new_n946), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n941), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n440), .B1(new_n708), .B2(new_n734), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n644), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n865), .B1(new_n932), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n932), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n223), .A2(new_n212), .A3(new_n584), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n531), .B(KEYINPUT102), .Z(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT35), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n961), .B1(new_n960), .B2(new_n959), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT36), .Z(new_n963));
  NOR3_X1   g0763(.A1(new_n705), .A2(new_n203), .A3(new_n331), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n229), .A2(G50), .ZN(new_n965));
  OAI211_X1 g0765(.A(G1), .B(new_n268), .C1(new_n964), .C2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n956), .A2(new_n963), .A3(new_n966), .ZN(G367));
  INV_X1    g0767(.A(KEYINPUT112), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n573), .A2(new_n671), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT110), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n970), .A2(new_n656), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n648), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n973), .A2(KEYINPUT111), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n973), .A2(KEYINPUT111), .ZN(new_n975));
  NOR3_X1   g0775(.A1(new_n974), .A2(new_n975), .A3(KEYINPUT43), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n714), .B(new_n721), .C1(new_n713), .C2(new_n672), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n651), .A2(new_n671), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(KEYINPUT42), .B1(new_n695), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n599), .A2(new_n672), .ZN(new_n982));
  AND2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n695), .A2(new_n697), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n697), .A2(KEYINPUT42), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n984), .A2(new_n979), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n973), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n976), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  INV_X1    g0790(.A(new_n976), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n983), .B2(new_n986), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n968), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n992), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n983), .A2(new_n986), .B1(KEYINPUT43), .B2(new_n988), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n994), .B(KEYINPUT112), .C1(new_n976), .C2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n693), .A2(new_n980), .ZN(new_n997));
  AND3_X1   g0797(.A1(new_n993), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n997), .B1(new_n993), .B2(new_n996), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n701), .B(KEYINPUT41), .Z(new_n1001));
  OAI21_X1  g0801(.A(new_n979), .B1(new_n698), .B2(new_n699), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT45), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(KEYINPUT45), .B(new_n979), .C1(new_n698), .C2(new_n699), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n984), .A2(KEYINPUT96), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n1008), .A3(new_n980), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT44), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1007), .A2(KEYINPUT44), .A3(new_n1008), .A4(new_n980), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1006), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n693), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1006), .A2(new_n1013), .A3(new_n693), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n695), .A2(KEYINPUT113), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n690), .B(new_n694), .C1(new_n686), .C2(new_n688), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n695), .A2(KEYINPUT113), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1021), .A2(new_n676), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(new_n676), .ZN(new_n1023));
  AND3_X1   g0823(.A1(new_n1022), .A2(new_n755), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1016), .A2(new_n1017), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1001), .B1(new_n1025), .B2(new_n755), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n758), .B(KEYINPUT114), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1000), .B1(new_n1026), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT46), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n794), .B2(new_n584), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n768), .B1(KEYINPUT115), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(KEYINPUT115), .B2(new_n1031), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n786), .A2(new_n604), .B1(new_n780), .B2(new_n829), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(G317), .B2(new_n809), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n789), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n793), .A2(G311), .B1(new_n1036), .B2(G97), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G107), .A2(new_n799), .B1(new_n800), .B2(G294), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n795), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n793), .A2(G143), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n229), .B2(new_n798), .C1(new_n203), .C2(new_n789), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n800), .A2(G159), .B1(new_n795), .B2(G58), .ZN(new_n1043));
  XOR2_X1   g0843(.A(KEYINPUT116), .B(G137), .Z(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n809), .A2(new_n1045), .B1(new_n815), .B2(G50), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n428), .B1(new_n787), .B2(G150), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1043), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n1033), .A2(new_n1040), .B1(new_n1042), .B2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT47), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n774), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n769), .A2(new_n252), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n776), .B1(new_n216), .B2(new_n565), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n759), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1051), .B(new_n1054), .C1(new_n988), .C2(new_n822), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1029), .A2(new_n1055), .ZN(G387));
  NOR2_X1   g0856(.A1(new_n692), .A2(new_n822), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(new_n787), .A2(G317), .B1(new_n815), .B2(G303), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n793), .A2(G322), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(new_n781), .C2(new_n806), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT48), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n799), .A2(G283), .B1(new_n795), .B2(G294), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT49), .ZN(new_n1066));
  OR2_X1    g0866(.A1(new_n1066), .A2(KEYINPUT118), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(KEYINPUT118), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n789), .A2(new_n584), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n1069), .B(new_n768), .C1(G326), .C2(new_n809), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n806), .A2(new_n276), .B1(new_n420), .B2(new_n798), .ZN(new_n1072));
  INV_X1    g0872(.A(G159), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n808), .A2(new_n1073), .B1(new_n794), .B2(new_n203), .ZN(new_n1074));
  NOR2_X1   g0874(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n786), .A2(new_n202), .B1(new_n780), .B2(new_n229), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(G150), .B2(new_n809), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n790), .A2(G97), .ZN(new_n1078));
  NAND4_X1  g0878(.A1(new_n1075), .A2(new_n768), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n826), .B1(new_n1071), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n418), .A2(new_n202), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT50), .Z(new_n1082));
  AOI21_X1  g0882(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1082), .A2(new_n703), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n249), .A2(G45), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n1084), .A2(new_n1085), .A3(new_n769), .ZN(new_n1086));
  OAI221_X1 g0886(.A(new_n1086), .B1(G107), .B2(new_n215), .C1(new_n703), .C2(new_n763), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n759), .B1(new_n1087), .B2(new_n775), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT117), .Z(new_n1089));
  NOR3_X1   g0889(.A1(new_n1057), .A2(new_n1080), .A3(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(new_n1021), .B(new_n675), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1090), .B1(new_n1091), .B2(new_n1028), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1091), .A2(new_n755), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n701), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1091), .A2(new_n755), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1092), .B1(new_n1094), .B2(new_n1095), .ZN(G393));
  AND3_X1   g0896(.A1(new_n1006), .A2(new_n1013), .A3(new_n693), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n693), .B1(new_n1006), .B2(new_n1013), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1093), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1099), .A2(new_n1025), .A3(new_n701), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n832), .A2(new_n841), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n418), .A2(new_n815), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n800), .A2(G50), .B1(G143), .B2(new_n809), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n798), .A2(new_n203), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n233), .B2(new_n795), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .A4(new_n1105), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G150), .A2(new_n793), .B1(new_n787), .B2(G159), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT51), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G317), .A2(new_n793), .B1(new_n787), .B2(G311), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT52), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n428), .B1(new_n780), .B2(new_n468), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(G322), .B2(new_n809), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n800), .A2(G303), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n799), .A2(G116), .B1(new_n795), .B2(G283), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n813), .A2(new_n1112), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1106), .A2(new_n1108), .B1(new_n1110), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n774), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n769), .A2(new_n256), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n1118), .B(new_n775), .C1(new_n206), .C2(new_n215), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n760), .A3(new_n1119), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1120), .B1(new_n980), .B2(new_n773), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1121), .B1(new_n1122), .B2(new_n1028), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1100), .A2(new_n1123), .ZN(G390));
  NAND4_X1  g0924(.A1(new_n904), .A2(new_n908), .A3(new_n909), .A4(G330), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n938), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(new_n934), .A2(new_n935), .B1(new_n947), .B2(new_n1127), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n898), .A2(new_n918), .A3(KEYINPUT108), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n938), .A2(KEYINPUT119), .ZN(new_n1130));
  INV_X1    g0930(.A(KEYINPUT119), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n936), .A2(new_n1131), .A3(new_n937), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1130), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n849), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n732), .B2(new_n848), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n946), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1133), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT108), .B1(new_n898), .B2(new_n918), .ZN(new_n1138));
  NOR3_X1   g0938(.A1(new_n1129), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1126), .B1(new_n1128), .B2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n1134), .B1(new_n856), .B2(new_n857), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1127), .B1(new_n1141), .B2(new_n1136), .ZN(new_n1142));
  AND3_X1   g0942(.A1(new_n891), .A2(KEYINPUT39), .A3(new_n898), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1142), .B1(new_n1143), .B2(new_n933), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n850), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n754), .A2(new_n1145), .A3(new_n946), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1137), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1147), .A2(new_n921), .A3(new_n922), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1144), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n440), .A2(new_n904), .A3(G330), .A4(new_n909), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n952), .A2(new_n644), .A3(new_n1150), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n904), .A2(new_n909), .A3(G330), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1136), .B1(new_n1152), .B2(new_n850), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1153), .A2(new_n1146), .A3(new_n1135), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n946), .B1(new_n754), .B2(new_n1145), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n945), .B1(new_n1126), .B2(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1151), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1140), .A2(new_n1149), .A3(new_n1157), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1157), .B(KEYINPUT120), .ZN(new_n1159));
  AND2_X1   g0959(.A1(new_n1140), .A2(new_n1149), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n701), .B(new_n1158), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1140), .A2(new_n1149), .A3(new_n1028), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n771), .B1(new_n1143), .B2(new_n933), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n760), .B1(new_n367), .B2(new_n827), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n806), .A2(new_n207), .B1(new_n808), .B2(new_n829), .ZN(new_n1165));
  AOI211_X1 g0965(.A(new_n1104), .B(new_n1165), .C1(G87), .C2(new_n795), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n786), .A2(new_n584), .B1(new_n780), .B2(new_n206), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n296), .B(new_n1167), .C1(G294), .C2(new_n809), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1166), .B(new_n1168), .C1(new_n229), .C2(new_n831), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT121), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n806), .A2(new_n1044), .B1(new_n789), .B2(new_n202), .ZN(new_n1171));
  INV_X1    g0971(.A(G128), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n808), .A2(new_n1172), .B1(new_n1073), .B2(new_n798), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT54), .B(G143), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n296), .B1(new_n780), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(G132), .ZN(new_n1177));
  INV_X1    g0977(.A(G125), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n786), .A2(new_n1177), .B1(new_n783), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n795), .A2(G150), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1176), .B(new_n1179), .C1(KEYINPUT53), .C2(new_n1180), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1174), .B(new_n1181), .C1(KEYINPUT53), .C2(new_n1180), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT122), .B1(new_n1170), .B2(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1183), .A2(new_n826), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1170), .A2(KEYINPUT122), .A3(new_n1182), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1164), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1163), .A2(new_n1186), .ZN(new_n1187));
  AND3_X1   g0987(.A1(new_n1162), .A2(KEYINPUT123), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(KEYINPUT123), .B1(new_n1162), .B2(new_n1187), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1161), .B1(new_n1188), .B2(new_n1189), .ZN(G378));
  NAND2_X1  g0990(.A1(new_n281), .A2(new_n871), .ZN(new_n1191));
  XNOR2_X1  g0991(.A(new_n313), .B(new_n1191), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1192), .B(new_n1193), .Z(new_n1194));
  AOI21_X1  g0994(.A(new_n910), .B1(new_n891), .B2(new_n898), .ZN(new_n1195));
  OAI21_X1  g0995(.A(G330), .B1(new_n1195), .B2(KEYINPUT40), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n1129), .A2(new_n1138), .A3(new_n923), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1194), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1192), .B(new_n1193), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n911), .A2(G330), .A3(new_n925), .A4(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1198), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n951), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1198), .A2(new_n1200), .A3(new_n941), .A4(new_n950), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n1028), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1194), .A2(new_n771), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n760), .B1(G50), .B2(new_n827), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n786), .A2(new_n1172), .B1(new_n780), .B2(new_n837), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1175), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n800), .A2(G132), .B1(new_n795), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n1178), .B2(new_n808), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1208), .B(new_n1211), .C1(G150), .C2(new_n799), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1036), .A2(G159), .ZN(new_n1216));
  AOI211_X1 g1016(.A(G33), .B(G41), .C1(new_n809), .C2(G124), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n841), .A2(new_n445), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n789), .A2(new_n330), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(G97), .B2(new_n800), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n584), .B2(new_n808), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n787), .A2(G107), .B1(new_n815), .B2(new_n565), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n829), .B2(new_n783), .ZN(new_n1224));
  OAI22_X1  g1024(.A1(new_n798), .A2(new_n229), .B1(new_n794), .B2(new_n203), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1219), .A2(new_n1222), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(KEYINPUT58), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1219), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1228));
  OR2_X1    g1028(.A1(new_n1226), .A2(KEYINPUT58), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1218), .A2(new_n1227), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1207), .B1(new_n1230), .B2(new_n774), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1206), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1205), .A2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1151), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n1202), .A2(new_n1203), .B1(new_n1234), .B2(new_n1158), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n702), .B1(new_n1235), .B2(KEYINPUT57), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1158), .A2(new_n1234), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1204), .A2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT57), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1233), .B1(new_n1236), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(G375));
  OAI21_X1  g1042(.A(new_n760), .B1(G68), .B2(new_n827), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n786), .A2(new_n829), .B1(new_n780), .B2(new_n207), .ZN(new_n1244));
  AOI211_X1 g1044(.A(new_n296), .B(new_n1244), .C1(G303), .C2(new_n809), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n790), .A2(G77), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n565), .A2(new_n799), .B1(new_n800), .B2(G116), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n793), .A2(G294), .B1(new_n795), .B2(G97), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1245), .A2(new_n1246), .A3(new_n1247), .A4(new_n1248), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n787), .A2(new_n1045), .B1(new_n815), .B2(G150), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1172), .B2(new_n783), .ZN(new_n1251));
  AOI211_X1 g1051(.A(new_n1220), .B(new_n1251), .C1(G132), .C2(new_n793), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n800), .A2(new_n1209), .B1(new_n795), .B2(G159), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1252), .B(new_n1253), .C1(new_n202), .C2(new_n798), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1249), .B1(new_n1254), .B2(new_n841), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1243), .B1(new_n1255), .B2(new_n774), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n946), .B2(new_n772), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1258), .B2(new_n1027), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1258), .A2(new_n1151), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1001), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1260), .B1(new_n1159), .B2(new_n1263), .ZN(G381));
  NOR4_X1   g1064(.A1(G381), .A2(G393), .A3(G396), .A4(G384), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1162), .A2(new_n1187), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1161), .A2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(G390), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1265), .A2(new_n1268), .A3(new_n1269), .ZN(new_n1270));
  OR3_X1    g1070(.A1(G375), .A2(G387), .A3(new_n1270), .ZN(G407));
  NAND2_X1  g1071(.A1(new_n670), .A2(G213), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1241), .A2(new_n1268), .A3(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(G407), .A2(G213), .A3(new_n1274), .ZN(G409));
  XNOR2_X1  g1075(.A(G393), .B(new_n824), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AND3_X1   g1077(.A1(new_n1029), .A2(new_n1055), .A3(G390), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G390), .B1(new_n1029), .B2(new_n1055), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1277), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n993), .A2(new_n996), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n997), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n993), .A2(new_n996), .A3(new_n997), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(new_n1097), .A2(new_n1098), .A3(new_n1093), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n755), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1262), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1285), .B1(new_n1288), .B2(new_n1027), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1055), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1269), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1029), .A2(new_n1055), .A3(G390), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1276), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1280), .A2(new_n1293), .ZN(new_n1294));
  INV_X1    g1094(.A(KEYINPUT60), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1261), .B1(new_n1157), .B2(new_n1295), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1258), .A2(KEYINPUT60), .A3(new_n1151), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1296), .A2(new_n701), .A3(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1298), .A2(new_n1260), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n863), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1298), .A2(G384), .A3(new_n1260), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1273), .A2(G2897), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(KEYINPUT126), .ZN(new_n1303));
  AND3_X1   g1103(.A1(new_n1300), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1304), .A2(new_n1305), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1201), .A2(new_n951), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n1198), .A2(new_n1200), .B1(new_n941), .B2(new_n950), .ZN(new_n1308));
  OAI211_X1 g1108(.A(new_n1237), .B(new_n1262), .C1(new_n1307), .C2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT124), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  AOI22_X1  g1111(.A1(new_n1204), .A2(new_n1028), .B1(new_n1206), .B2(new_n1231), .ZN(new_n1312));
  NAND4_X1  g1112(.A1(new_n1204), .A2(KEYINPUT124), .A3(new_n1262), .A4(new_n1237), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1311), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  AOI22_X1  g1114(.A1(new_n1241), .A2(G378), .B1(new_n1314), .B2(new_n1268), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1306), .B1(new_n1315), .B2(new_n1273), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1314), .A2(new_n1268), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1204), .A2(KEYINPUT57), .A3(new_n1237), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n701), .ZN(new_n1319));
  NOR2_X1   g1119(.A1(new_n1235), .A2(KEYINPUT57), .ZN(new_n1320));
  OAI211_X1 g1120(.A(G378), .B(new_n1312), .C1(new_n1319), .C2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1317), .A2(new_n1321), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT62), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1322), .A2(new_n1323), .A3(new_n1272), .A4(new_n1324), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT61), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1316), .A2(new_n1325), .A3(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1273), .B1(new_n1317), .B2(new_n1321), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1323), .B1(new_n1328), .B2(new_n1324), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1294), .B1(new_n1327), .B2(new_n1329), .ZN(new_n1330));
  AOI211_X1 g1130(.A(KEYINPUT125), .B(KEYINPUT63), .C1(new_n1328), .C2(new_n1324), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT125), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1322), .A2(new_n1272), .A3(new_n1324), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT63), .ZN(new_n1334));
  AOI21_X1  g1134(.A(new_n1332), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1331), .A2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(new_n1280), .A2(new_n1326), .A3(new_n1293), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1337), .A2(KEYINPUT127), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1328), .A2(KEYINPUT63), .A3(new_n1324), .ZN(new_n1339));
  INV_X1    g1139(.A(KEYINPUT127), .ZN(new_n1340));
  NAND4_X1  g1140(.A1(new_n1280), .A2(new_n1293), .A3(new_n1340), .A4(new_n1326), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1338), .A2(new_n1316), .A3(new_n1339), .A4(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1330), .B1(new_n1336), .B2(new_n1342), .ZN(G405));
  OAI21_X1  g1143(.A(new_n1321), .B1(new_n1241), .B2(new_n1267), .ZN(new_n1344));
  XNOR2_X1  g1144(.A(new_n1344), .B(new_n1324), .ZN(new_n1345));
  XNOR2_X1  g1145(.A(new_n1345), .B(new_n1294), .ZN(G402));
endmodule


