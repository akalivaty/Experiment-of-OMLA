//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0005(.A(G50), .B1(G58), .B2(G68), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NAND2_X1  g0007(.A1(G1), .A2(G13), .ZN(new_n208));
  NOR3_X1   g0008(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT0), .ZN(new_n213));
  AOI21_X1  g0013(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G116), .ZN(new_n218));
  INV_X1    g0018(.A(G270), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n210), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n214), .B1(new_n213), .B2(new_n212), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G226), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT64), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n231), .B(new_n235), .Z(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  XNOR2_X1  g0043(.A(KEYINPUT3), .B(G33), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n244), .A2(G223), .A3(G1698), .ZN(new_n245));
  INV_X1    g0045(.A(G77), .ZN(new_n246));
  INV_X1    g0046(.A(G1698), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G222), .ZN(new_n249));
  OAI221_X1 g0049(.A(new_n245), .B1(new_n246), .B2(new_n244), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(G33), .A2(G41), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n251), .A2(G1), .A3(G13), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  AND2_X1   g0054(.A1(G33), .A2(G41), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G41), .A2(G45), .ZN(new_n256));
  OAI22_X1  g0056(.A1(new_n255), .A2(new_n208), .B1(new_n256), .B2(G1), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT66), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT66), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n260), .B1(G41), .B2(G45), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n252), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G226), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT65), .B(G45), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n260), .B(G274), .C1(new_n265), .C2(G41), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n254), .A2(new_n264), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G190), .ZN(new_n268));
  OR2_X1    g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(G200), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G20), .A2(G33), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n207), .A2(G33), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT8), .B(G58), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n208), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n202), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n277), .B1(new_n260), .B2(G20), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n280), .B1(new_n281), .B2(new_n202), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(new_n283), .B(KEYINPUT9), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n269), .A2(new_n270), .A3(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(new_n285), .B(KEYINPUT10), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n267), .A2(G169), .ZN(new_n287));
  INV_X1    g0087(.A(G179), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n287), .B1(new_n288), .B2(new_n267), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n283), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT17), .ZN(new_n292));
  INV_X1    g0092(.A(new_n274), .ZN(new_n293));
  INV_X1    g0093(.A(new_n279), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n281), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n295), .B1(new_n296), .B2(new_n293), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT7), .ZN(new_n299));
  NOR3_X1   g0099(.A1(new_n244), .A2(new_n299), .A3(G20), .ZN(new_n300));
  INV_X1    g0100(.A(G33), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT3), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT3), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G33), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g0105(.A(KEYINPUT7), .B1(new_n305), .B2(new_n207), .ZN(new_n306));
  OAI21_X1  g0106(.A(G68), .B1(new_n300), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G58), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(new_n216), .ZN(new_n309));
  OAI21_X1  g0109(.A(G20), .B1(new_n309), .B2(new_n201), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n271), .A2(G159), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n307), .A2(KEYINPUT16), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n277), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n299), .A2(G20), .ZN(new_n316));
  OAI21_X1  g0116(.A(KEYINPUT72), .B1(new_n303), .B2(G33), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n304), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n302), .A2(KEYINPUT72), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n316), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n299), .B1(new_n244), .B2(G20), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G68), .ZN(new_n323));
  AOI21_X1  g0123(.A(KEYINPUT16), .B1(new_n323), .B2(new_n313), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n298), .B1(new_n315), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n252), .A2(G232), .A3(new_n261), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n266), .A2(new_n326), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n302), .A2(new_n304), .A3(G226), .A4(G1698), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT73), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT73), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n244), .A2(new_n330), .A3(G226), .A4(G1698), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G87), .ZN(new_n332));
  NAND4_X1  g0132(.A1(new_n302), .A2(new_n304), .A3(G223), .A4(new_n247), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n329), .A2(new_n331), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  AOI211_X1 g0134(.A(G190), .B(new_n327), .C1(new_n334), .C2(new_n253), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n332), .B(new_n333), .C1(new_n328), .C2(KEYINPUT73), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n328), .A2(KEYINPUT73), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n253), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n327), .ZN(new_n339));
  AOI21_X1  g0139(.A(G200), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n335), .A2(new_n340), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n292), .B1(new_n325), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n277), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n305), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n321), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n312), .B1(new_n345), .B2(G68), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n343), .B1(new_n346), .B2(KEYINPUT16), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT16), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n216), .B1(new_n320), .B2(new_n321), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n348), .B1(new_n349), .B2(new_n312), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n297), .B1(new_n347), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n338), .A2(new_n288), .A3(new_n339), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n327), .B1(new_n334), .B2(new_n253), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(G169), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT18), .B1(new_n351), .B2(new_n354), .ZN(new_n355));
  AOI211_X1 g0155(.A(G179), .B(new_n327), .C1(new_n334), .C2(new_n253), .ZN(new_n356));
  AOI21_X1  g0156(.A(G169), .B1(new_n338), .B2(new_n339), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT18), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n325), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n338), .A2(new_n268), .A3(new_n339), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(G200), .B2(new_n353), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n351), .A2(KEYINPUT17), .A3(new_n362), .ZN(new_n363));
  NAND4_X1  g0163(.A1(new_n342), .A2(new_n355), .A3(new_n360), .A4(new_n363), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT15), .B(G87), .ZN(new_n365));
  OR2_X1    g0165(.A1(new_n365), .A2(new_n273), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT68), .B1(new_n207), .B2(new_n246), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT68), .ZN(new_n369));
  XOR2_X1   g0169(.A(new_n274), .B(KEYINPUT67), .Z(new_n370));
  INV_X1    g0170(.A(new_n271), .ZN(new_n371));
  OAI221_X1 g0171(.A(new_n368), .B1(new_n369), .B2(new_n366), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n277), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n279), .A2(new_n246), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n281), .B2(new_n246), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n305), .A2(G107), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n244), .A2(G1698), .ZN(new_n378));
  OAI221_X1 g0178(.A(new_n377), .B1(new_n248), .B2(new_n230), .C1(new_n217), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n253), .ZN(new_n380));
  INV_X1    g0180(.A(new_n266), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n381), .B1(G244), .B2(new_n263), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n380), .A2(new_n382), .A3(new_n268), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n380), .A2(new_n382), .ZN(new_n384));
  INV_X1    g0184(.A(G200), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n376), .B1(new_n383), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(G169), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n288), .B2(new_n384), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n376), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NOR4_X1   g0191(.A1(new_n291), .A2(new_n364), .A3(new_n387), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n260), .A2(G13), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(G20), .A3(new_n216), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT12), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n216), .B2(new_n296), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n371), .A2(new_n202), .B1(new_n207), .B2(G68), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n273), .A2(new_n246), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n277), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT11), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n400), .A2(new_n401), .ZN(new_n404));
  NOR3_X1   g0204(.A1(new_n397), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  AND3_X1   g0206(.A1(new_n252), .A2(new_n259), .A3(new_n261), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n259), .B1(new_n252), .B2(new_n261), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n407), .A2(new_n408), .A3(KEYINPUT69), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT69), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n410), .B1(new_n258), .B2(new_n262), .ZN(new_n411));
  OAI21_X1  g0211(.A(G238), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT70), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(new_n266), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT69), .B1(new_n407), .B2(new_n408), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n258), .A2(new_n410), .A3(new_n262), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n217), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT70), .B1(new_n417), .B2(new_n381), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n244), .A2(G226), .A3(new_n247), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G97), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n419), .B(new_n420), .C1(new_n378), .C2(new_n230), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(new_n253), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n414), .A2(new_n418), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT13), .ZN(new_n424));
  INV_X1    g0224(.A(new_n422), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n415), .A2(new_n416), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n381), .B1(new_n426), .B2(G238), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n425), .B1(new_n427), .B2(new_n413), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT13), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(new_n418), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n424), .A2(new_n430), .A3(G179), .ZN(new_n431));
  INV_X1    g0231(.A(G169), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n424), .B2(new_n430), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT14), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n431), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  AOI211_X1 g0235(.A(KEYINPUT14), .B(new_n432), .C1(new_n424), .C2(new_n430), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n406), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n424), .A2(new_n430), .A3(G190), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n405), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT71), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n424), .A2(new_n430), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n442), .B2(G200), .ZN(new_n443));
  AOI211_X1 g0243(.A(KEYINPUT71), .B(new_n385), .C1(new_n424), .C2(new_n430), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n440), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AND3_X1   g0245(.A1(new_n392), .A2(new_n437), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT75), .ZN(new_n447));
  XNOR2_X1  g0247(.A(KEYINPUT5), .B(G41), .ZN(new_n448));
  INV_X1    g0248(.A(G45), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(G1), .ZN(new_n450));
  INV_X1    g0250(.A(new_n208), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n448), .A2(new_n450), .B1(new_n451), .B2(new_n251), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n447), .B1(new_n452), .B2(G257), .ZN(new_n453));
  INV_X1    g0253(.A(G41), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT5), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT5), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(G41), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n450), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND4_X1  g0258(.A1(new_n458), .A2(new_n447), .A3(G257), .A4(new_n252), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n448), .A2(G274), .A3(new_n450), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g0261(.A(KEYINPUT76), .B1(new_n453), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(G33), .A2(G283), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n302), .A2(new_n304), .A3(G244), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT4), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n244), .A2(KEYINPUT4), .A3(G244), .A4(new_n247), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n466), .B1(new_n244), .B2(G250), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n467), .B(new_n468), .C1(new_n247), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n253), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n458), .A2(G257), .A3(new_n252), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(KEYINPUT75), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT76), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n473), .A2(new_n474), .A3(new_n459), .A4(new_n460), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n462), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n385), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n477), .B1(G190), .B2(new_n476), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n294), .A2(G97), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n260), .A2(G33), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n279), .A2(new_n480), .A3(new_n208), .A4(new_n276), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n479), .B1(G97), .B2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT74), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT6), .ZN(new_n484));
  INV_X1    g0284(.A(G97), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n484), .A2(new_n485), .A3(G107), .ZN(new_n486));
  XNOR2_X1  g0286(.A(G97), .B(G107), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n486), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  OAI221_X1 g0288(.A(new_n483), .B1(new_n246), .B2(new_n371), .C1(new_n488), .C2(new_n207), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n487), .A2(new_n484), .ZN(new_n490));
  INV_X1    g0290(.A(new_n486), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n207), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n371), .A2(new_n246), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT74), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n322), .A2(G107), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n489), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n482), .B1(new_n496), .B2(new_n277), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n478), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n462), .A2(new_n471), .A3(new_n288), .A4(new_n475), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT77), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n473), .A2(new_n459), .A3(new_n460), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n501), .A2(KEYINPUT76), .B1(new_n470), .B2(new_n253), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT77), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n502), .A2(new_n503), .A3(new_n288), .A4(new_n475), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n496), .A2(new_n277), .ZN(new_n506));
  INV_X1    g0306(.A(new_n482), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n506), .A2(new_n507), .B1(new_n476), .B2(new_n432), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n498), .A2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n207), .A2(G107), .ZN(new_n512));
  AOI21_X1  g0312(.A(KEYINPUT25), .B1(new_n394), .B2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT83), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G107), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n515), .B1(new_n516), .B2(new_n481), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n394), .A2(new_n512), .A3(KEYINPUT25), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT83), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n519), .A2(new_n513), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT82), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n302), .A2(new_n304), .A3(new_n207), .A4(G87), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT22), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT22), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n244), .A2(new_n526), .A3(new_n207), .A4(G87), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT23), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n529), .A2(new_n516), .A3(G20), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n531));
  OAI21_X1  g0331(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n530), .B(new_n531), .C1(new_n532), .C2(KEYINPUT81), .ZN(new_n533));
  AND2_X1   g0333(.A1(new_n532), .A2(KEYINPUT81), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n528), .A2(new_n535), .A3(KEYINPUT24), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n277), .ZN(new_n537));
  AOI21_X1  g0337(.A(KEYINPUT24), .B1(new_n528), .B2(new_n535), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n523), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n528), .A2(new_n535), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT24), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n542), .A2(KEYINPUT82), .A3(new_n277), .A4(new_n536), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n522), .B1(new_n539), .B2(new_n543), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n302), .A2(new_n304), .A3(G257), .A4(G1698), .ZN(new_n545));
  INV_X1    g0345(.A(G294), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n301), .B2(new_n546), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n244), .A2(G250), .A3(new_n247), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n253), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n458), .A2(G264), .A3(new_n252), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(KEYINPUT84), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT84), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n452), .A2(new_n552), .A3(G264), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n549), .A2(new_n460), .A3(new_n551), .A4(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(new_n288), .ZN(new_n555));
  AND2_X1   g0355(.A1(new_n550), .A2(new_n460), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n432), .B1(new_n549), .B2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n544), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n549), .A2(new_n268), .A3(new_n556), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n554), .A2(new_n385), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n544), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(G274), .ZN(new_n566));
  NOR2_X1   g0366(.A1(new_n458), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n567), .B1(G270), .B2(new_n452), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n302), .A2(new_n304), .A3(G264), .A4(G1698), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n302), .A2(new_n304), .A3(G257), .A4(new_n247), .ZN(new_n570));
  INV_X1    g0370(.A(G303), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n244), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n253), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n568), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n385), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n575), .B1(G190), .B2(new_n574), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n301), .A2(G97), .ZN(new_n577));
  AOI21_X1  g0377(.A(G20), .B1(new_n577), .B2(new_n463), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n207), .A2(new_n218), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n277), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT20), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(KEYINPUT20), .B(new_n277), .C1(new_n578), .C2(new_n579), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n481), .A2(G116), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(G116), .B2(new_n294), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n576), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(new_n586), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(KEYINPUT80), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n588), .A2(G169), .A3(new_n574), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n458), .A2(new_n252), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n460), .B1(new_n592), .B2(new_n219), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n253), .B2(new_n572), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n588), .A2(G179), .A3(new_n594), .ZN(new_n595));
  AND2_X1   g0395(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n588), .A2(G169), .A3(new_n574), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n597), .A2(KEYINPUT80), .A3(new_n589), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n587), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n365), .A2(new_n294), .ZN(new_n600));
  OR2_X1    g0400(.A1(new_n481), .A2(new_n365), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT19), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n207), .B1(new_n420), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(G87), .A2(G97), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n516), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n302), .A2(new_n304), .A3(new_n207), .A4(G68), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n207), .A2(G33), .A3(G97), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n602), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n606), .A2(new_n607), .A3(KEYINPUT78), .A4(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(new_n277), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n603), .A2(new_n605), .B1(new_n602), .B2(new_n608), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT78), .B1(new_n612), .B2(new_n607), .ZN(new_n613));
  OAI211_X1 g0413(.A(new_n600), .B(new_n601), .C1(new_n611), .C2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(G250), .B1(new_n449), .B2(G1), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n260), .A2(G45), .A3(G274), .ZN(new_n616));
  AOI22_X1  g0416(.A1(new_n615), .A2(new_n616), .B1(new_n451), .B2(new_n251), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n302), .A2(new_n304), .A3(G238), .A4(new_n247), .ZN(new_n618));
  NAND2_X1  g0418(.A1(G33), .A2(G116), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n618), .B(new_n619), .C1(new_n465), .C2(new_n247), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n617), .B1(new_n620), .B2(new_n253), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n288), .ZN(new_n622));
  AND2_X1   g0422(.A1(new_n614), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n621), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(new_n432), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n621), .A2(new_n385), .ZN(new_n626));
  AOI211_X1 g0426(.A(new_n268), .B(new_n617), .C1(new_n620), .C2(new_n253), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n600), .B1(new_n611), .B2(new_n613), .ZN(new_n629));
  INV_X1    g0429(.A(G87), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n481), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g0431(.A(new_n631), .B(KEYINPUT79), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n623), .A2(new_n625), .B1(new_n628), .B2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n599), .A2(new_n635), .ZN(new_n636));
  AND4_X1   g0436(.A1(new_n446), .A2(new_n511), .A3(new_n565), .A4(new_n636), .ZN(G372));
  AOI21_X1  g0437(.A(new_n429), .B1(new_n428), .B2(new_n418), .ZN(new_n638));
  AND4_X1   g0438(.A1(new_n429), .A2(new_n414), .A3(new_n418), .A4(new_n422), .ZN(new_n639));
  OAI21_X1  g0439(.A(G169), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(KEYINPUT14), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n442), .A2(new_n434), .A3(G169), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n641), .A2(new_n642), .A3(new_n431), .ZN(new_n643));
  AOI22_X1  g0443(.A1(new_n445), .A2(new_n391), .B1(new_n643), .B2(new_n406), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n342), .A2(new_n363), .ZN(new_n645));
  OAI211_X1 g0445(.A(new_n355), .B(new_n360), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n646), .A2(new_n286), .B1(new_n283), .B2(new_n289), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT85), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n620), .A2(new_n648), .A3(new_n253), .ZN(new_n649));
  INV_X1    g0449(.A(new_n617), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n648), .B1(new_n620), .B2(new_n253), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n432), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n623), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n596), .B(new_n598), .C1(new_n544), .C2(new_n558), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n657), .A2(new_n509), .A3(new_n498), .A4(new_n563), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n649), .A2(new_n650), .ZN(new_n659));
  OAI21_X1  g0459(.A(G200), .B1(new_n659), .B2(new_n652), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n633), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(KEYINPUT86), .ZN(new_n662));
  INV_X1    g0462(.A(new_n627), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT86), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n660), .A2(new_n633), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n662), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n656), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n656), .B1(new_n658), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n634), .A2(new_n505), .A3(new_n508), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT26), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n666), .A2(new_n505), .A3(new_n508), .A4(new_n656), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(KEYINPUT26), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n446), .B1(new_n668), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n647), .A2(new_n673), .ZN(G369));
  OR3_X1    g0474(.A1(new_n393), .A2(KEYINPUT27), .A3(G20), .ZN(new_n675));
  OAI21_X1  g0475(.A(KEYINPUT27), .B1(new_n393), .B2(G20), .ZN(new_n676));
  AND3_X1   g0476(.A1(new_n675), .A2(G213), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(G343), .ZN(new_n678));
  XOR2_X1   g0478(.A(new_n678), .B(KEYINPUT87), .Z(new_n679));
  NAND3_X1  g0479(.A1(new_n657), .A2(new_n563), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(G330), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n679), .B1(new_n584), .B2(new_n586), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT88), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n682), .B1(new_n599), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n683), .B2(new_n599), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n598), .A2(new_n591), .A3(new_n595), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n681), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  XOR2_X1   g0488(.A(new_n688), .B(KEYINPUT89), .Z(new_n689));
  NOR2_X1   g0489(.A1(new_n544), .A2(new_n679), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n564), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n679), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n559), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n680), .B1(new_n689), .B2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n211), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n604), .A2(new_n516), .A3(new_n218), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n700), .A2(G1), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n703), .B1(new_n206), .B2(new_n700), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT28), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n679), .B1(new_n668), .B2(new_n672), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT93), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT29), .ZN(new_n709));
  OAI211_X1 g0509(.A(KEYINPUT93), .B(new_n679), .C1(new_n668), .C2(new_n672), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n708), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n668), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT26), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n669), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT94), .ZN(new_n715));
  INV_X1    g0515(.A(new_n509), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(KEYINPUT26), .A3(new_n656), .A4(new_n666), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT94), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n669), .A2(new_n718), .A3(new_n713), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n715), .A2(new_n717), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n693), .B1(new_n712), .B2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT29), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n711), .A2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT31), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n679), .A2(new_n724), .ZN(new_n725));
  XOR2_X1   g0525(.A(KEYINPUT90), .B(KEYINPUT30), .Z(new_n726));
  AND3_X1   g0526(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(G179), .A3(new_n594), .A4(new_n621), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n726), .B1(new_n728), .B2(new_n476), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT91), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n594), .A2(G179), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n654), .A2(new_n476), .A3(new_n731), .A4(new_n554), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n729), .A2(new_n730), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n549), .A2(new_n551), .A3(new_n553), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n568), .A2(new_n573), .A3(G179), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n734), .A2(new_n735), .A3(new_n624), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(KEYINPUT30), .A3(new_n475), .A4(new_n502), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n733), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n730), .B1(new_n729), .B2(new_n732), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n725), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT92), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n729), .A2(new_n737), .A3(new_n732), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n693), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(new_n724), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n740), .A2(new_n741), .A3(new_n744), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n565), .A2(new_n511), .A3(new_n636), .A4(new_n679), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n741), .B1(new_n740), .B2(new_n744), .ZN(new_n748));
  OAI21_X1  g0548(.A(G330), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n723), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n705), .B1(new_n751), .B2(G1), .ZN(G364));
  NAND3_X1  g0552(.A1(new_n207), .A2(G13), .A3(G45), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n700), .A2(G1), .A3(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n685), .A2(new_n681), .A3(new_n687), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n755), .B1(new_n689), .B2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G13), .A2(G33), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G20), .ZN(new_n760));
  AND3_X1   g0560(.A1(new_n685), .A2(new_n687), .A3(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n208), .B1(G20), .B2(new_n432), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n698), .A2(new_n244), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n766), .B1(new_n206), .B2(new_n265), .C1(new_n239), .C2(new_n449), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n698), .A2(new_n305), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n768), .A2(G355), .B1(new_n218), .B2(new_n698), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n765), .B1(new_n767), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n207), .A2(G190), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G179), .A2(G200), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n773), .A2(KEYINPUT96), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(KEYINPUT96), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n771), .A2(new_n288), .A3(G200), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT97), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT97), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n777), .A2(G329), .B1(new_n782), .B2(G283), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n207), .A2(new_n268), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n288), .A2(new_n385), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n244), .B1(new_n787), .B2(G326), .ZN(new_n788));
  INV_X1    g0588(.A(new_n784), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n789), .A2(new_n385), .A3(G179), .ZN(new_n790));
  INV_X1    g0590(.A(new_n771), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n791), .A2(new_n288), .A3(G200), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G303), .A2(new_n790), .B1(new_n792), .B2(G311), .ZN(new_n793));
  NOR3_X1   g0593(.A1(new_n789), .A2(new_n288), .A3(G200), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G322), .ZN(new_n795));
  XOR2_X1   g0595(.A(KEYINPUT33), .B(G317), .Z(new_n796));
  NAND2_X1  g0596(.A1(new_n785), .A2(new_n771), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AND4_X1   g0598(.A1(new_n788), .A2(new_n793), .A3(new_n795), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n207), .B1(new_n772), .B2(G190), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n800), .A2(KEYINPUT99), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(KEYINPUT99), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n783), .B(new_n799), .C1(new_n546), .C2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n777), .A2(G159), .ZN(new_n805));
  INV_X1    g0605(.A(KEYINPUT32), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n803), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G97), .ZN(new_n809));
  INV_X1    g0609(.A(new_n792), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n810), .A2(new_n246), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n786), .A2(new_n202), .B1(new_n797), .B2(new_n216), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n794), .B(KEYINPUT95), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n811), .B(new_n812), .C1(new_n814), .C2(G58), .ZN(new_n815));
  AND3_X1   g0615(.A1(new_n807), .A2(new_n809), .A3(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n782), .A2(G107), .ZN(new_n818));
  INV_X1    g0618(.A(new_n790), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n818), .B(new_n244), .C1(new_n630), .C2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT98), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n804), .B1(new_n817), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n770), .B1(new_n822), .B2(new_n763), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n754), .B1(new_n762), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n757), .A2(new_n824), .ZN(G396));
  OAI22_X1  g0625(.A1(new_n819), .A2(new_n516), .B1(new_n810), .B2(new_n218), .ZN(new_n826));
  INV_X1    g0626(.A(new_n794), .ZN(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n827), .A2(new_n546), .B1(new_n797), .B2(new_n828), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n305), .B1(new_n786), .B2(new_n571), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n826), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n782), .A2(G87), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n777), .A2(G311), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n831), .A2(new_n809), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  AOI22_X1  g0634(.A1(new_n792), .A2(G159), .B1(new_n787), .B2(G137), .ZN(new_n835));
  INV_X1    g0635(.A(G150), .ZN(new_n836));
  INV_X1    g0636(.A(G143), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n835), .B1(new_n836), .B2(new_n797), .C1(new_n813), .C2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT34), .Z(new_n839));
  NOR2_X1   g0639(.A1(new_n781), .A2(new_n216), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n305), .B(new_n840), .C1(G50), .C2(new_n790), .ZN(new_n841));
  INV_X1    g0641(.A(G132), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n841), .B1(new_n308), .B2(new_n803), .C1(new_n842), .C2(new_n776), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n834), .B1(new_n839), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n763), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n763), .A2(new_n758), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n754), .B1(new_n246), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n391), .A2(new_n679), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n679), .B1(new_n373), .B2(new_n375), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n390), .B1(new_n387), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n845), .B(new_n847), .C1(new_n852), .C2(new_n759), .ZN(new_n853));
  INV_X1    g0653(.A(KEYINPUT100), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n708), .A2(new_n710), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n854), .B1(new_n855), .B2(new_n851), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n708), .A2(new_n854), .A3(new_n710), .A4(new_n851), .ZN(new_n857));
  OAI211_X1 g0657(.A(new_n679), .B(new_n852), .C1(new_n668), .C2(new_n672), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  OR3_X1    g0659(.A1(new_n856), .A2(new_n749), .A3(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT101), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n861), .B(new_n749), .C1(new_n856), .C2(new_n859), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n754), .A3(new_n862), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n856), .A2(new_n859), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n861), .B1(new_n864), .B2(new_n749), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n853), .B1(new_n863), .B2(new_n865), .ZN(G384));
  AOI21_X1  g0666(.A(new_n260), .B1(G13), .B2(new_n207), .ZN(new_n867));
  OAI21_X1  g0667(.A(G200), .B1(new_n638), .B2(new_n639), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT71), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n442), .A2(new_n441), .A3(G200), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n439), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI211_X1 g0671(.A(new_n406), .B(new_n693), .C1(new_n871), .C2(new_n643), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n693), .A2(new_n406), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n437), .A2(new_n445), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n743), .B(KEYINPUT31), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n746), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT38), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT37), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n216), .B1(new_n321), .B2(new_n344), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n348), .B1(new_n880), .B2(new_n312), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n314), .A2(new_n881), .A3(new_n277), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n298), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT102), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n882), .A2(KEYINPUT102), .A3(new_n298), .ZN(new_n886));
  INV_X1    g0686(.A(new_n677), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n354), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n885), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n351), .A2(new_n362), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n879), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n325), .A2(new_n358), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n325), .A2(new_n677), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n892), .A2(new_n893), .A3(new_n890), .A4(new_n879), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n882), .A2(KEYINPUT102), .A3(new_n298), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT102), .B1(new_n882), .B2(new_n298), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n897), .A2(new_n898), .A3(new_n887), .ZN(new_n899));
  AND2_X1   g0699(.A1(new_n364), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n878), .B1(new_n896), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n364), .A2(new_n899), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n902), .B(KEYINPUT38), .C1(new_n895), .C2(new_n891), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n875), .A2(new_n852), .A3(new_n877), .A4(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT40), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n851), .B1(new_n872), .B2(new_n874), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n892), .A2(new_n893), .A3(new_n890), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  INV_X1    g0710(.A(new_n893), .ZN(new_n911));
  AOI22_X1  g0711(.A1(new_n910), .A2(new_n894), .B1(new_n364), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n912), .A2(KEYINPUT38), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n906), .B1(new_n914), .B2(new_n903), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n908), .A2(new_n915), .A3(new_n877), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n907), .A2(new_n916), .ZN(new_n917));
  XOR2_X1   g0717(.A(new_n917), .B(KEYINPUT105), .Z(new_n918));
  AND2_X1   g0718(.A1(new_n446), .A2(new_n877), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n681), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n918), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n711), .A2(new_n446), .A3(new_n722), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT104), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND4_X1  g0724(.A1(new_n711), .A2(new_n446), .A3(KEYINPUT104), .A4(new_n722), .ZN(new_n925));
  AND3_X1   g0725(.A1(new_n924), .A2(new_n647), .A3(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n643), .A2(new_n406), .A3(new_n679), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT39), .ZN(new_n929));
  OAI211_X1 g0729(.A(new_n903), .B(new_n929), .C1(KEYINPUT38), .C2(new_n912), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n929), .B1(new_n901), .B2(new_n903), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n858), .A2(new_n848), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n875), .A3(new_n904), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n355), .A2(new_n360), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n887), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n933), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT103), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT103), .ZN(new_n940));
  NAND4_X1  g0740(.A1(new_n933), .A2(new_n935), .A3(new_n940), .A4(new_n937), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n926), .B(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n867), .B1(new_n921), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n921), .B2(new_n943), .ZN(new_n945));
  NOR3_X1   g0745(.A1(new_n309), .A2(new_n206), .A3(new_n246), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n202), .B2(G68), .ZN(new_n947));
  OR3_X1    g0747(.A1(new_n947), .A2(new_n260), .A3(G13), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n208), .A2(new_n207), .A3(new_n218), .ZN(new_n949));
  INV_X1    g0749(.A(new_n488), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n949), .B1(new_n950), .B2(KEYINPUT35), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(KEYINPUT35), .B2(new_n950), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT36), .Z(new_n953));
  NAND3_X1  g0753(.A1(new_n945), .A2(new_n948), .A3(new_n953), .ZN(G367));
  INV_X1    g0754(.A(new_n763), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n819), .A2(new_n308), .B1(new_n810), .B2(new_n202), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n244), .B1(new_n827), .B2(new_n836), .ZN(new_n957));
  INV_X1    g0757(.A(G159), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n786), .A2(new_n837), .B1(new_n797), .B2(new_n958), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n956), .A2(new_n957), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n808), .A2(G68), .ZN(new_n961));
  XOR2_X1   g0761(.A(KEYINPUT112), .B(G137), .Z(new_n962));
  NAND2_X1  g0762(.A1(new_n777), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n782), .A2(G77), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n960), .A2(new_n961), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n790), .A2(G116), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT46), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n808), .A2(G107), .ZN(new_n968));
  INV_X1    g0768(.A(new_n797), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n244), .B1(new_n969), .B2(G294), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n792), .A2(G283), .B1(new_n787), .B2(G311), .ZN(new_n971));
  NAND4_X1  g0771(.A1(new_n967), .A2(new_n968), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n777), .A2(G317), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n782), .A2(G97), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n973), .B(new_n974), .C1(new_n571), .C2(new_n813), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n965), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n955), .B1(new_n977), .B2(KEYINPUT47), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(KEYINPUT47), .B2(new_n977), .ZN(new_n979));
  INV_X1    g0779(.A(new_n766), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n235), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n764), .B1(new_n211), .B2(new_n365), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n979), .B(new_n755), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n983), .B(KEYINPUT113), .ZN(new_n984));
  INV_X1    g0784(.A(new_n760), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n679), .A2(new_n633), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(new_n656), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT106), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n666), .A2(new_n656), .A3(new_n986), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n984), .B1(new_n985), .B2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n679), .A2(new_n497), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n510), .A2(new_n992), .B1(new_n509), .B2(new_n679), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n693), .B1(new_n596), .B2(new_n598), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n691), .A2(new_n993), .A3(new_n994), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT42), .Z(new_n996));
  AOI21_X1  g0796(.A(new_n716), .B1(new_n498), .B2(new_n559), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n996), .B1(new_n693), .B2(new_n997), .ZN(new_n998));
  INV_X1    g0798(.A(KEYINPUT107), .ZN(new_n999));
  OR2_X1    g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n998), .A2(new_n999), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n990), .A2(KEYINPUT43), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g0805(.A(new_n990), .B(KEYINPUT43), .Z(new_n1006));
  INV_X1    g0806(.A(new_n1006), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1000), .A2(new_n1007), .A3(new_n1001), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n689), .A2(new_n696), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n993), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(KEYINPUT108), .ZN(new_n1014));
  INV_X1    g0814(.A(KEYINPUT108), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1009), .A2(new_n1015), .A3(new_n1012), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1005), .A2(new_n1011), .A3(new_n1008), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1014), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n753), .A2(G1), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n993), .A2(new_n680), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT45), .Z(new_n1021));
  NOR2_X1   g0821(.A1(new_n993), .A2(new_n680), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT44), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  AND3_X1   g0824(.A1(new_n1010), .A2(KEYINPUT109), .A3(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(KEYINPUT109), .B1(new_n1010), .B2(new_n1024), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1010), .A2(new_n1024), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n691), .A2(new_n994), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(new_n695), .B2(new_n994), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n689), .A2(new_n1031), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT111), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n689), .A2(new_n1031), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT110), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1034), .B(new_n1035), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n751), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n699), .B(KEYINPUT41), .Z(new_n1039));
  INV_X1    g0839(.A(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1019), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n991), .B1(new_n1018), .B2(new_n1041), .ZN(G387));
  NOR2_X1   g0842(.A1(new_n1037), .A2(new_n750), .ZN(new_n1043));
  INV_X1    g0843(.A(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1037), .A2(new_n750), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(new_n699), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1037), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(KEYINPUT115), .B(G322), .ZN(new_n1048));
  AOI22_X1  g0848(.A1(new_n787), .A2(new_n1048), .B1(new_n969), .B2(G311), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n571), .B2(new_n810), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1050), .B1(new_n814), .B2(G317), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT48), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(KEYINPUT48), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n808), .A2(G283), .B1(G294), .B2(new_n790), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT49), .ZN(new_n1056));
  OR2_X1    g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n305), .B1(new_n781), .B2(new_n218), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(G326), .B2(new_n777), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1057), .A2(new_n1058), .A3(new_n1060), .ZN(new_n1061));
  OAI22_X1  g0861(.A1(new_n810), .A2(new_n216), .B1(new_n274), .B2(new_n797), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n819), .A2(new_n246), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n827), .A2(new_n202), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n244), .B1(new_n786), .B2(new_n958), .ZN(new_n1065));
  NOR4_X1   g0865(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .A4(new_n1065), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n803), .A2(new_n365), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n777), .A2(G150), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n1066), .A2(new_n974), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n955), .B1(new_n1061), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n231), .A2(new_n265), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n370), .A2(G50), .ZN(new_n1073));
  XOR2_X1   g0873(.A(KEYINPUT114), .B(KEYINPUT50), .Z(new_n1074));
  XNOR2_X1  g0874(.A(new_n1073), .B(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n702), .B(new_n449), .C1(new_n216), .C2(new_n246), .ZN(new_n1076));
  OAI211_X1 g0876(.A(new_n1072), .B(new_n766), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n768), .A2(new_n701), .B1(new_n516), .B2(new_n698), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n765), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NOR3_X1   g0879(.A1(new_n1071), .A2(new_n754), .A3(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT116), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n696), .A2(new_n760), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1047), .A2(new_n1019), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1046), .A2(new_n1083), .ZN(G393));
  INV_X1    g0884(.A(new_n1027), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1010), .A2(new_n1024), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n1086), .A3(new_n1019), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n764), .B1(new_n485), .B2(new_n211), .C1(new_n242), .C2(new_n980), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n755), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n244), .B1(new_n202), .B2(new_n797), .C1(new_n819), .C2(new_n216), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G87), .B2(new_n782), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n1091), .B1(new_n837), .B2(new_n776), .C1(new_n370), .C2(new_n810), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n794), .A2(G159), .B1(new_n787), .B2(G150), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n803), .A2(new_n246), .ZN(new_n1095));
  OR2_X1    g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n777), .A2(new_n1048), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n244), .B1(new_n792), .B2(G294), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n790), .A2(G283), .B1(G303), .B2(new_n969), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1097), .A2(new_n818), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n794), .A2(G311), .B1(new_n787), .B2(G317), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT52), .Z(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n218), .B2(new_n803), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n1092), .A2(new_n1096), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1089), .B1(new_n1104), .B2(new_n763), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n993), .B2(new_n985), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1087), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1044), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n700), .B1(new_n1043), .B2(new_n1028), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1107), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(G390));
  INV_X1    g0912(.A(new_n875), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n681), .B1(new_n876), .B2(new_n746), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1114), .A2(KEYINPUT117), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n852), .B1(new_n1114), .B2(KEYINPUT117), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1113), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n715), .A2(new_n717), .A3(new_n719), .ZN(new_n1118));
  OAI211_X1 g0918(.A(new_n679), .B(new_n850), .C1(new_n1118), .C2(new_n668), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n848), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n749), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n1120), .B1(new_n1121), .B2(new_n908), .ZN(new_n1122));
  OAI211_X1 g0922(.A(G330), .B(new_n852), .C1(new_n747), .C2(new_n748), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1113), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n908), .A2(new_n1114), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1117), .A2(new_n1122), .B1(new_n1126), .B2(new_n934), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n446), .A2(G330), .A3(new_n877), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n924), .A2(new_n647), .A3(new_n925), .A4(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1125), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n903), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n325), .A2(new_n341), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n897), .A2(new_n898), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(new_n1135), .B2(new_n888), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n894), .B1(new_n1136), .B2(new_n879), .ZN(new_n1137));
  AOI21_X1  g0937(.A(KEYINPUT38), .B1(new_n1137), .B2(new_n902), .ZN(new_n1138));
  OAI21_X1  g0938(.A(KEYINPUT39), .B1(new_n1133), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n930), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n934), .A2(new_n875), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n927), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n927), .B1(new_n1133), .B2(new_n913), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1143), .B1(new_n1120), .B2(new_n875), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1132), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1143), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n848), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1147), .B1(new_n721), .B2(new_n850), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1146), .B1(new_n1148), .B2(new_n1113), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n931), .A2(new_n932), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n848), .A2(new_n858), .B1(new_n872), .B2(new_n874), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n928), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1121), .A2(new_n908), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1149), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1145), .A2(new_n1154), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1131), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1155), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n699), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1145), .A2(new_n1154), .A3(new_n1019), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n846), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n755), .B1(new_n293), .B2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(G128), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n244), .B1(new_n786), .B2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n827), .A2(new_n842), .ZN(new_n1164));
  AOI211_X1 g0964(.A(new_n1163), .B(new_n1164), .C1(new_n969), .C2(new_n962), .ZN(new_n1165));
  OAI221_X1 g0965(.A(new_n1165), .B1(new_n202), .B2(new_n781), .C1(new_n958), .C2(new_n803), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n790), .A2(G150), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT53), .Z(new_n1168));
  XNOR2_X1  g0968(.A(KEYINPUT54), .B(G143), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT118), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(new_n792), .ZN(new_n1171));
  INV_X1    g0971(.A(G125), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1168), .B(new_n1171), .C1(new_n1172), .C2(new_n776), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n840), .B1(G294), .B2(new_n777), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n244), .B1(new_n790), .B2(G87), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n794), .A2(G116), .B1(new_n787), .B2(G283), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n792), .A2(G97), .B1(new_n969), .B2(G107), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1174), .A2(new_n1175), .A3(new_n1176), .A4(new_n1177), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n1166), .A2(new_n1173), .B1(new_n1095), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1161), .B1(new_n1179), .B2(new_n763), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1180), .B1(new_n1140), .B2(new_n759), .ZN(new_n1181));
  AND3_X1   g0981(.A1(new_n1159), .A2(KEYINPUT119), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT119), .B1(new_n1159), .B2(new_n1181), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n1156), .A2(new_n1158), .B1(new_n1182), .B2(new_n1183), .ZN(G378));
  NAND3_X1  g0984(.A1(new_n939), .A2(KEYINPUT122), .A3(new_n941), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n907), .A2(G330), .A3(new_n916), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n283), .A2(new_n677), .ZN(new_n1187));
  XNOR2_X1  g0987(.A(new_n291), .B(new_n1187), .ZN(new_n1188));
  XOR2_X1   g0988(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1189));
  XNOR2_X1  g0989(.A(new_n1188), .B(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1186), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1190), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1192), .A2(new_n907), .A3(G330), .A4(new_n916), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n1185), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1185), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1190), .A2(new_n758), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n755), .B1(G50), .B2(new_n1160), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n786), .A2(new_n1172), .B1(new_n797), .B2(new_n842), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G137), .B2(new_n792), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1170), .A2(new_n790), .B1(G128), .B2(new_n794), .ZN(new_n1201));
  AND2_X1   g1001(.A1(new_n1201), .A2(KEYINPUT120), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1201), .A2(KEYINPUT120), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1200), .B1(new_n836), .B2(new_n803), .C1(new_n1202), .C2(new_n1203), .ZN(new_n1204));
  XOR2_X1   g1004(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1205));
  OR2_X1    g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n301), .B(new_n454), .C1(new_n781), .C2(new_n958), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(G124), .B2(new_n777), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1209), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n827), .A2(new_n516), .B1(new_n797), .B2(new_n485), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n810), .A2(new_n365), .B1(new_n218), .B2(new_n786), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n305), .A2(new_n454), .ZN(new_n1213));
  NOR4_X1   g1013(.A1(new_n1211), .A2(new_n1212), .A3(new_n1063), .A4(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n782), .A2(G58), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n777), .A2(G283), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1214), .A2(new_n961), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT58), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1213), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1210), .A2(new_n1219), .A3(new_n1220), .A4(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1198), .B1(new_n1222), .B2(new_n763), .ZN(new_n1223));
  AOI22_X1  g1023(.A1(new_n1196), .A2(new_n1019), .B1(new_n1197), .B2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n926), .B(new_n1128), .C1(new_n1155), .C2(new_n1127), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n942), .A2(new_n1191), .A3(new_n1193), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n942), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1225), .B(KEYINPUT57), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT123), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1228), .A2(new_n1229), .A3(new_n699), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1225), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT57), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1230), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1229), .B1(new_n1228), .B2(new_n699), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1224), .B1(new_n1234), .B2(new_n1235), .ZN(G375));
  NAND2_X1  g1036(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1131), .A2(new_n1040), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1113), .A2(new_n758), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n755), .B1(G68), .B2(new_n1160), .ZN(new_n1240));
  OAI22_X1  g1040(.A1(new_n810), .A2(new_n836), .B1(new_n842), .B2(new_n786), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n305), .B(new_n1241), .C1(G159), .C2(new_n790), .ZN(new_n1242));
  OAI211_X1 g1042(.A(new_n1242), .B(new_n1215), .C1(new_n202), .C2(new_n803), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n814), .A2(new_n962), .B1(new_n969), .B2(new_n1170), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n1162), .B2(new_n776), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n485), .A2(new_n819), .B1(new_n827), .B2(new_n828), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n810), .A2(new_n516), .B1(new_n797), .B2(new_n218), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n244), .B1(new_n787), .B2(G294), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n777), .A2(G303), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1248), .A2(new_n964), .A3(new_n1249), .A4(new_n1250), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n1243), .A2(new_n1245), .B1(new_n1067), .B2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1240), .B1(new_n1252), .B2(new_n763), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1239), .A2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1019), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1254), .B1(new_n1127), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1238), .A2(new_n1257), .ZN(G381));
  OAI211_X1 g1058(.A(new_n1046), .B(new_n1083), .C1(new_n757), .C2(new_n824), .ZN(new_n1259));
  OR2_X1    g1059(.A1(new_n1259), .A2(G384), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n750), .B1(new_n1047), .B2(new_n1028), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1255), .B1(new_n1261), .B2(new_n1039), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1262), .A2(new_n1014), .A3(new_n1016), .A4(new_n1017), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(new_n991), .A3(new_n1111), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1159), .A2(new_n1181), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1224), .B(new_n1267), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1268));
  OR4_X1    g1068(.A1(G381), .A2(new_n1260), .A3(new_n1264), .A4(new_n1268), .ZN(G407));
  OAI211_X1 g1069(.A(G407), .B(G213), .C1(G343), .C2(new_n1268), .ZN(G409));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  INV_X1    g1071(.A(G343), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(G213), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  OAI211_X1 g1074(.A(G378), .B(new_n1224), .C1(new_n1234), .C2(new_n1235), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1197), .A2(new_n1223), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1019), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1276), .B(new_n1277), .C1(new_n1231), .C2(new_n1039), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1267), .A2(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1274), .B1(new_n1275), .B2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1274), .A2(G2897), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(G384), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT124), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n699), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1237), .A2(KEYINPUT60), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT60), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1127), .A2(new_n1129), .A3(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1285), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1283), .B(new_n1284), .C1(new_n1289), .C2(new_n1256), .ZN(new_n1290));
  AND3_X1   g1090(.A1(new_n1127), .A2(new_n1129), .A3(new_n1287), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1287), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  OAI211_X1 g1093(.A(G384), .B(new_n1257), .C1(new_n1293), .C2(new_n1285), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1290), .A2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1257), .B1(new_n1293), .B2(new_n1285), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1284), .B1(new_n1296), .B2(new_n1283), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1282), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1283), .B1(new_n1289), .B2(new_n1256), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT124), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1300), .A2(new_n1290), .A3(new_n1294), .A4(new_n1281), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1298), .A2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1271), .B1(new_n1280), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(KEYINPUT126), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT126), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1305), .B(new_n1271), .C1(new_n1280), .C2(new_n1302), .ZN(new_n1306));
  NOR2_X1   g1106(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1280), .A2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1308), .A2(KEYINPUT62), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1280), .A2(new_n1310), .A3(new_n1307), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1304), .A2(new_n1306), .A3(new_n1309), .A4(new_n1311), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(G393), .A2(G396), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1259), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  NOR2_X1   g1115(.A1(G387), .A2(G390), .ZN(new_n1316));
  AOI21_X1  g1116(.A(new_n1111), .B1(new_n1263), .B2(new_n991), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1315), .B1(new_n1316), .B2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(G387), .A2(G390), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1319), .A2(new_n1264), .A3(new_n1314), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1312), .A2(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1321), .A2(KEYINPUT61), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1280), .A2(KEYINPUT63), .A3(new_n1307), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1280), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1298), .A2(KEYINPUT125), .A3(new_n1301), .ZN(new_n1326));
  AOI21_X1  g1126(.A(KEYINPUT125), .B1(new_n1298), .B2(new_n1301), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1325), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT63), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1308), .A2(new_n1329), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1323), .A2(new_n1324), .A3(new_n1328), .A4(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1322), .A2(new_n1331), .ZN(G405));
  INV_X1    g1132(.A(KEYINPUT127), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(G375), .A2(new_n1267), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(new_n1275), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1335), .A2(new_n1307), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1307), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1334), .A2(new_n1337), .A3(new_n1275), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1321), .A2(new_n1333), .A3(new_n1336), .A4(new_n1338), .ZN(new_n1339));
  AND2_X1   g1139(.A1(new_n1336), .A2(new_n1338), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1339), .B1(new_n1321), .B2(new_n1340), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1333), .B1(new_n1340), .B2(new_n1321), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1341), .A2(new_n1342), .ZN(G402));
endmodule


