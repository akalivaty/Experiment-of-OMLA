//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n847, new_n848, new_n850,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n972, new_n973, new_n974,
    new_n975, new_n976;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  OAI21_X1  g002(.A(KEYINPUT92), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n202), .A2(new_n203), .A3(KEYINPUT14), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT14), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT92), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n208), .A2(G29gat), .A3(G36gat), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n204), .A2(new_n205), .A3(new_n207), .A4(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT15), .ZN(new_n211));
  XOR2_X1   g010(.A(G43gat), .B(G50gat), .Z(new_n212));
  AOI21_X1  g011(.A(new_n211), .B1(new_n212), .B2(KEYINPUT89), .ZN(new_n213));
  XNOR2_X1  g012(.A(G43gat), .B(G50gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT89), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(new_n210), .B1(new_n213), .B2(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(KEYINPUT90), .B(G43gat), .Z(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(G50gat), .ZN(new_n219));
  XOR2_X1   g018(.A(KEYINPUT91), .B(G50gat), .Z(new_n220));
  NOR2_X1   g019(.A1(new_n220), .A2(G43gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n211), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n217), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(KEYINPUT15), .B1(new_n214), .B2(new_n215), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n224), .B1(new_n215), .B2(new_n214), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n205), .B(new_n207), .C1(new_n202), .C2(new_n203), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT17), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n231), .A2(G1gat), .ZN(new_n232));
  INV_X1    g031(.A(G8gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n231), .B1(new_n234), .B2(G1gat), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n233), .B1(new_n232), .B2(new_n235), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI22_X1  g037(.A1(new_n222), .A2(new_n217), .B1(new_n225), .B2(new_n226), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT17), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n230), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G229gat), .A2(G233gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n238), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n241), .A2(KEYINPUT18), .A3(new_n242), .A4(new_n244), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n238), .B1(new_n239), .B2(KEYINPUT17), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n223), .A2(KEYINPUT17), .A3(new_n227), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n242), .B(new_n244), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT18), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n239), .A2(new_n238), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n244), .A2(new_n251), .ZN(new_n252));
  XOR2_X1   g051(.A(new_n242), .B(KEYINPUT13), .Z(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G113gat), .B(G141gat), .ZN(new_n255));
  XNOR2_X1  g054(.A(G169gat), .B(G197gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT12), .ZN(new_n260));
  AND4_X1   g059(.A1(new_n245), .A2(new_n250), .A3(new_n254), .A4(new_n260), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n248), .A2(new_n249), .B1(new_n252), .B2(new_n253), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n260), .B1(new_n262), .B2(new_n245), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT93), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n261), .A2(new_n263), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT93), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(G113gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT72), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(G113gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n273), .A3(G120gat), .ZN(new_n274));
  OR3_X1    g073(.A1(new_n270), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT71), .B1(new_n270), .B2(G120gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  OR2_X1    g076(.A1(G127gat), .A2(G134gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(G127gat), .A2(G134gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(KEYINPUT1), .B1(new_n280), .B2(KEYINPUT73), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(new_n282), .A3(new_n279), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n277), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT2), .ZN(new_n285));
  INV_X1    g084(.A(G141gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(G148gat), .ZN(new_n287));
  INV_X1    g086(.A(G148gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(G141gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n285), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G155gat), .ZN(new_n291));
  INV_X1    g090(.A(G162gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G155gat), .A2(G162gat), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT81), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n296), .B1(new_n286), .B2(G148gat), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n288), .A2(KEYINPUT81), .A3(G141gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n286), .A2(G148gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n294), .B1(new_n293), .B2(KEYINPUT2), .ZN(new_n301));
  AOI22_X1  g100(.A1(new_n290), .A2(new_n295), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G134gat), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n303), .A2(KEYINPUT70), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n303), .A2(KEYINPUT70), .ZN(new_n305));
  OAI21_X1  g104(.A(G127gat), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT1), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n270), .A2(G120gat), .ZN(new_n308));
  INV_X1    g107(.A(G120gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(G113gat), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n307), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n306), .A2(new_n311), .A3(new_n278), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n284), .A2(new_n302), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT4), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n284), .A2(new_n302), .A3(new_n315), .A4(new_n312), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n290), .A2(new_n295), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n300), .A2(new_n301), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT82), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT82), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(KEYINPUT3), .A3(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT3), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n312), .A2(new_n284), .B1(new_n302), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  AND2_X1   g126(.A1(new_n317), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G225gat), .A2(G233gat), .ZN(new_n329));
  NOR3_X1   g128(.A1(new_n328), .A2(KEYINPUT39), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G1gat), .B(G29gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(KEYINPUT0), .ZN(new_n332));
  XNOR2_X1  g131(.A(G57gat), .B(G85gat), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n332), .B(new_n333), .Z(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  AND3_X1   g135(.A1(new_n274), .A2(new_n276), .A3(new_n275), .ZN(new_n337));
  INV_X1    g136(.A(new_n279), .ZN(new_n338));
  NOR2_X1   g137(.A1(G127gat), .A2(G134gat), .ZN(new_n339));
  OAI21_X1  g138(.A(KEYINPUT73), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(new_n283), .A3(new_n307), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n312), .B1(new_n337), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n321), .A2(new_n342), .A3(new_n323), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n343), .A2(new_n329), .A3(new_n313), .ZN(new_n344));
  OAI211_X1 g143(.A(KEYINPUT39), .B(new_n344), .C1(new_n328), .C2(new_n329), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n336), .A2(KEYINPUT40), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT40), .B1(new_n336), .B2(new_n345), .ZN(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n343), .A2(new_n313), .ZN(new_n349));
  INV_X1    g148(.A(new_n329), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n317), .A2(new_n327), .A3(new_n329), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n317), .A2(new_n327), .A3(new_n329), .A4(new_n348), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n334), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n346), .A2(new_n347), .A3(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G8gat), .B(G36gat), .Z(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(KEYINPUT80), .ZN(new_n358));
  XNOR2_X1  g157(.A(G64gat), .B(G92gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n358), .B(new_n359), .Z(new_n360));
  INV_X1    g159(.A(G169gat), .ZN(new_n361));
  INV_X1    g160(.A(G176gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT23), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT23), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n364), .B1(G169gat), .B2(G176gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(G169gat), .A2(G176gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n368), .B1(G183gat), .B2(G190gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(G183gat), .A2(G190gat), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT24), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT64), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(KEYINPUT64), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n367), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT65), .B1(new_n376), .B2(KEYINPUT25), .ZN(new_n377));
  INV_X1    g176(.A(G183gat), .ZN(new_n378));
  INV_X1    g177(.A(G190gat), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n370), .B1(KEYINPUT67), .B2(KEYINPUT24), .ZN(new_n381));
  AND2_X1   g180(.A1(KEYINPUT67), .A2(KEYINPUT24), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n380), .B(new_n368), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n365), .A2(KEYINPUT25), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n363), .A2(KEYINPUT66), .A3(new_n366), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT66), .B1(new_n363), .B2(new_n366), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n383), .B(new_n384), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT68), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT65), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT25), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n374), .A2(KEYINPUT64), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n392), .A2(new_n369), .A3(new_n372), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n390), .B(new_n391), .C1(new_n393), .C2(new_n367), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n363), .A2(new_n366), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT66), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n363), .A2(KEYINPUT66), .A3(new_n366), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n399), .A2(KEYINPUT68), .A3(new_n383), .A4(new_n384), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n377), .A2(new_n389), .A3(new_n394), .A4(new_n400), .ZN(new_n401));
  NOR2_X1   g200(.A1(G169gat), .A2(G176gat), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n402), .A2(KEYINPUT26), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n366), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n402), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n405));
  OR2_X1    g204(.A1(new_n378), .A2(KEYINPUT69), .ZN(new_n406));
  AOI21_X1  g205(.A(G190gat), .B1(new_n406), .B2(KEYINPUT27), .ZN(new_n407));
  OR3_X1    g206(.A1(new_n378), .A2(KEYINPUT69), .A3(KEYINPUT27), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT28), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  XOR2_X1   g208(.A(KEYINPUT27), .B(G183gat), .Z(new_n410));
  INV_X1    g209(.A(KEYINPUT28), .ZN(new_n411));
  NOR3_X1   g210(.A1(new_n410), .A2(new_n411), .A3(G190gat), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n404), .B(new_n405), .C1(new_n409), .C2(new_n412), .ZN(new_n413));
  AND2_X1   g212(.A1(G226gat), .A2(G233gat), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n401), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n414), .A2(KEYINPUT29), .ZN(new_n417));
  INV_X1    g216(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n401), .B2(new_n413), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT79), .ZN(new_n420));
  XNOR2_X1  g219(.A(G211gat), .B(G218gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT78), .ZN(new_n422));
  XNOR2_X1  g221(.A(G197gat), .B(G204gat), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n423), .B1(new_n421), .B2(KEYINPUT78), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(KEYINPUT76), .B(KEYINPUT22), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT77), .ZN(new_n427));
  INV_X1    g226(.A(G218gat), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(KEYINPUT77), .A2(G218gat), .ZN(new_n430));
  AND2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(G211gat), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n426), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n422), .B1(new_n425), .B2(new_n433), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n432), .B1(new_n429), .B2(new_n430), .ZN(new_n435));
  XOR2_X1   g234(.A(KEYINPUT76), .B(KEYINPUT22), .Z(new_n436));
  NOR2_X1   g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n422), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n437), .A2(new_n438), .A3(new_n424), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n420), .B1(new_n434), .B2(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n425), .A2(new_n433), .A3(new_n422), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n438), .B1(new_n437), .B2(new_n424), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT79), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n440), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NOR3_X1   g244(.A1(new_n416), .A2(new_n419), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n401), .A2(new_n413), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n417), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n444), .B1(new_n448), .B2(new_n415), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n360), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n445), .B1(new_n416), .B2(new_n419), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n448), .A2(new_n444), .A3(new_n415), .ZN(new_n452));
  INV_X1    g251(.A(new_n360), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n450), .A2(KEYINPUT30), .A3(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT30), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n451), .A2(new_n452), .A3(new_n456), .A4(new_n453), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n455), .A2(KEYINPUT87), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT87), .B1(new_n455), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n356), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G78gat), .B(G106gat), .ZN(new_n461));
  XNOR2_X1  g260(.A(KEYINPUT31), .B(G50gat), .ZN(new_n462));
  XOR2_X1   g261(.A(new_n461), .B(new_n462), .Z(new_n463));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G228gat), .A2(G233gat), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT29), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n441), .A2(new_n442), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(new_n325), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n321), .A2(new_n323), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n467), .B1(new_n320), .B2(KEYINPUT3), .ZN(new_n474));
  AOI22_X1  g273(.A1(new_n472), .A2(new_n473), .B1(new_n444), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n470), .B1(new_n325), .B2(new_n468), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT85), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n466), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n441), .A2(new_n442), .A3(KEYINPUT79), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT79), .B1(new_n441), .B2(new_n442), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n474), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n469), .A2(new_n320), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n481), .A2(new_n482), .A3(new_n466), .ZN(new_n483));
  NOR3_X1   g282(.A1(new_n478), .A2(new_n483), .A3(G22gat), .ZN(new_n484));
  INV_X1    g283(.A(G22gat), .ZN(new_n485));
  INV_X1    g284(.A(new_n466), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n481), .B1(new_n476), .B2(KEYINPUT85), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n472), .A2(new_n473), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n483), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n465), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(G22gat), .B1(new_n478), .B2(new_n483), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n489), .A2(new_n485), .A3(new_n490), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n463), .B(KEYINPUT86), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n493), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT37), .B1(new_n446), .B2(new_n449), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT37), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n451), .A2(new_n452), .A3(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n499), .A2(new_n360), .A3(new_n501), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n502), .A2(KEYINPUT38), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(KEYINPUT38), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n355), .A2(KEYINPUT6), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n353), .A2(new_n334), .A3(new_n354), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(new_n505), .B(new_n454), .C1(new_n508), .C2(new_n355), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n503), .A2(new_n504), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n460), .A2(new_n498), .A3(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(new_n342), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n447), .A2(new_n513), .ZN(new_n514));
  AND2_X1   g313(.A1(G227gat), .A2(G233gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n401), .A2(new_n342), .A3(new_n413), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(KEYINPUT32), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT33), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  XOR2_X1   g319(.A(G15gat), .B(G43gat), .Z(new_n521));
  XNOR2_X1  g320(.A(G71gat), .B(G99gat), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n518), .A2(new_n520), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n523), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n517), .B(KEYINPUT32), .C1(new_n519), .C2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT75), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n515), .B1(new_n514), .B2(new_n516), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT34), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n530), .B1(KEYINPUT74), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(KEYINPUT74), .B(KEYINPUT34), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n532), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n527), .A2(new_n528), .A3(new_n534), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n536), .A2(KEYINPUT36), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n535), .A2(new_n527), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT36), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n534), .A2(new_n524), .A3(new_n526), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n353), .A2(new_n354), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(new_n335), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT84), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n506), .A2(new_n507), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n355), .A2(KEYINPUT84), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AOI22_X1  g349(.A1(new_n550), .A2(new_n505), .B1(new_n457), .B2(new_n455), .ZN(new_n551));
  OR2_X1    g350(.A1(new_n551), .A2(new_n498), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n512), .A2(new_n543), .A3(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n551), .A2(new_n536), .A3(new_n537), .A4(new_n498), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n554), .A2(KEYINPUT35), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n458), .A2(new_n459), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n548), .A2(new_n545), .ZN(new_n558));
  AOI21_X1  g357(.A(KEYINPUT35), .B1(new_n558), .B2(new_n505), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n556), .A2(new_n557), .A3(new_n498), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n269), .B1(new_n553), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G71gat), .A2(G78gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(G71gat), .A2(G78gat), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(G57gat), .ZN(new_n566));
  INV_X1    g365(.A(G64gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g367(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n563), .B(new_n565), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(KEYINPUT94), .A2(G57gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(new_n567), .ZN(new_n572));
  INV_X1    g371(.A(new_n563), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(KEYINPUT9), .B2(new_n564), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n570), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(KEYINPUT95), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT95), .ZN(new_n577));
  OAI211_X1 g376(.A(new_n577), .B(new_n570), .C1(new_n572), .C2(new_n574), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n243), .B1(KEYINPUT21), .B2(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n579), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT21), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n586), .A2(G231gat), .A3(G233gat), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n586), .B1(G231gat), .B2(G233gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G127gat), .B(G155gat), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n590), .B(KEYINPUT96), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  XOR2_X1   g392(.A(G183gat), .B(G211gat), .Z(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n591), .B1(new_n587), .B2(new_n588), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n593), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n595), .B1(new_n593), .B2(new_n596), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n583), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n593), .A2(new_n596), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(new_n594), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n593), .A2(new_n596), .A3(new_n595), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n601), .A2(new_n582), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(G232gat), .A2(G233gat), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n605), .A2(KEYINPUT41), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT97), .ZN(new_n607));
  XOR2_X1   g406(.A(G134gat), .B(G162gat), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n609), .B(KEYINPUT100), .ZN(new_n610));
  XNOR2_X1  g409(.A(G99gat), .B(G106gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(G99gat), .ZN(new_n614));
  INV_X1    g413(.A(G106gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G99gat), .A2(G106gat), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n616), .A2(KEYINPUT98), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n613), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G85gat), .ZN(new_n620));
  INV_X1    g419(.A(G92gat), .ZN(new_n621));
  AOI22_X1  g420(.A1(KEYINPUT8), .A2(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT7), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n623), .B1(new_n620), .B2(new_n621), .ZN(new_n624));
  NAND3_X1  g423(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n619), .B(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n627), .B1(new_n228), .B2(new_n229), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n240), .ZN(new_n629));
  XNOR2_X1  g428(.A(G190gat), .B(G218gat), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT99), .Z(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n228), .A2(new_n627), .B1(KEYINPUT41), .B2(new_n605), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n632), .B1(new_n629), .B2(new_n633), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n610), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n629), .A2(new_n633), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n631), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n609), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n629), .A2(new_n632), .A3(new_n633), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n638), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n604), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT10), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n568), .A2(new_n569), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n573), .A2(new_n564), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n571), .B(G64gat), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT9), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n563), .B1(new_n565), .B2(new_n649), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n646), .A2(new_n647), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT101), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n626), .A2(new_n652), .A3(new_n613), .A4(new_n618), .ZN(new_n653));
  AND2_X1   g452(.A1(new_n624), .A2(new_n625), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT101), .B1(new_n654), .B2(new_n622), .ZN(new_n655));
  INV_X1    g454(.A(new_n619), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n651), .B(new_n653), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(new_n645), .B(new_n657), .C1(new_n579), .C2(new_n627), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT102), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n579), .A2(new_n627), .A3(KEYINPUT10), .ZN(new_n660));
  AND3_X1   g459(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n659), .B1(new_n658), .B2(new_n660), .ZN(new_n662));
  NAND2_X1  g461(.A1(G230gat), .A2(G233gat), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR3_X1   g463(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n657), .B1(new_n579), .B2(new_n627), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n664), .ZN(new_n667));
  XOR2_X1   g466(.A(G120gat), .B(G148gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n668), .B(KEYINPUT103), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n665), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n664), .B1(new_n658), .B2(new_n660), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n671), .B1(new_n675), .B2(new_n667), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n644), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n562), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n550), .A2(new_n505), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G1gat), .ZN(G1324gat));
  INV_X1    g484(.A(new_n556), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n233), .B1(new_n681), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT16), .B(G8gat), .ZN(new_n688));
  NOR3_X1   g487(.A1(new_n680), .A2(new_n556), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT42), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(KEYINPUT42), .B2(new_n689), .ZN(G1325gat));
  OAI21_X1  g490(.A(G15gat), .B1(new_n680), .B2(new_n543), .ZN(new_n692));
  INV_X1    g491(.A(new_n557), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(G15gat), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n692), .B1(new_n680), .B2(new_n694), .ZN(G1326gat));
  INV_X1    g494(.A(new_n498), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n697), .B(KEYINPUT104), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  INV_X1    g499(.A(new_n604), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n677), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n643), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n562), .A2(new_n703), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n704), .A2(G29gat), .A3(new_n682), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT45), .Z(new_n706));
  NOR2_X1   g505(.A1(new_n702), .A2(new_n267), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n553), .A2(new_n561), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT105), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n553), .A2(new_n561), .A3(KEYINPUT105), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n643), .A2(KEYINPUT44), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n643), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n709), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(KEYINPUT44), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n708), .B1(new_n714), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n682), .ZN(new_n720));
  AND2_X1   g519(.A1(new_n720), .A2(KEYINPUT106), .ZN(new_n721));
  OAI21_X1  g520(.A(G29gat), .B1(new_n720), .B2(KEYINPUT106), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n706), .B1(new_n721), .B2(new_n722), .ZN(G1328gat));
  NOR3_X1   g522(.A1(new_n704), .A2(G36gat), .A3(new_n556), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT46), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n719), .A2(new_n556), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n726), .A2(KEYINPUT107), .ZN(new_n727));
  OAI21_X1  g526(.A(G36gat), .B1(new_n726), .B2(KEYINPUT107), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(G1329gat));
  NAND2_X1  g528(.A1(new_n557), .A2(new_n218), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n704), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(KEYINPUT47), .B1(new_n732), .B2(KEYINPUT108), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT109), .ZN(new_n735));
  INV_X1    g534(.A(new_n543), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n718), .A2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(new_n218), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n735), .B1(new_n739), .B2(new_n732), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n218), .B1(new_n718), .B2(new_n736), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n741), .A2(KEYINPUT109), .A3(new_n731), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n734), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n739), .A2(new_n735), .A3(new_n732), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT109), .B1(new_n741), .B2(new_n731), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(new_n733), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(G1330gat));
  OAI21_X1  g546(.A(new_n220), .B1(new_n704), .B2(new_n498), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n498), .A2(new_n220), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n748), .B1(new_n719), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g550(.A1(new_n711), .A2(new_n712), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n644), .A2(new_n264), .A3(new_n677), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n682), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(new_n566), .ZN(G1332gat));
  NOR2_X1   g555(.A1(new_n754), .A2(new_n556), .ZN(new_n757));
  NOR2_X1   g556(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n758));
  AND2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n757), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n757), .B2(new_n758), .ZN(G1333gat));
  OAI21_X1  g560(.A(G71gat), .B1(new_n754), .B2(new_n543), .ZN(new_n762));
  INV_X1    g561(.A(G71gat), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n557), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n754), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g565(.A1(new_n754), .A2(new_n498), .ZN(new_n767));
  XOR2_X1   g566(.A(new_n767), .B(G78gat), .Z(G1335gat));
  NAND2_X1  g567(.A1(new_n714), .A2(new_n717), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n264), .A2(new_n677), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n769), .A2(new_n701), .A3(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(G85gat), .B1(new_n771), .B2(new_n682), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n604), .A2(new_n264), .ZN(new_n773));
  AND4_X1   g572(.A1(KEYINPUT51), .A2(new_n709), .A3(new_n715), .A4(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n643), .B1(new_n553), .B2(new_n561), .ZN(new_n775));
  AOI21_X1  g574(.A(KEYINPUT51), .B1(new_n775), .B2(new_n773), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n683), .A2(new_n620), .A3(new_n678), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT110), .Z(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n772), .A2(new_n780), .ZN(G1336gat));
  OAI21_X1  g580(.A(G92gat), .B1(new_n771), .B2(new_n556), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n556), .A2(G92gat), .A3(new_n677), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n784), .B2(KEYINPUT111), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n785), .B(new_n787), .ZN(G1337gat));
  OAI21_X1  g587(.A(G99gat), .B1(new_n771), .B2(new_n543), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n777), .A2(new_n614), .A3(new_n557), .A4(new_n678), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(G1338gat));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n498), .A2(G106gat), .A3(new_n677), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n774), .B2(new_n776), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n701), .A2(new_n770), .ZN(new_n795));
  AOI211_X1 g594(.A(new_n498), .B(new_n795), .C1(new_n714), .C2(new_n717), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n792), .B(new_n794), .C1(new_n796), .C2(new_n615), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(KEYINPUT112), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT112), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n799), .B(new_n793), .C1(new_n774), .C2(new_n776), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n798), .B(new_n800), .C1(new_n796), .C2(new_n615), .ZN(new_n801));
  AND3_X1   g600(.A1(new_n801), .A2(KEYINPUT113), .A3(KEYINPUT53), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT113), .B1(new_n801), .B2(KEYINPUT53), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n797), .B1(new_n802), .B2(new_n803), .ZN(G1339gat));
  NAND4_X1  g603(.A1(new_n604), .A2(new_n267), .A3(new_n643), .A4(new_n677), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT55), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n658), .A2(new_n664), .A3(new_n660), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT54), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n658), .A2(new_n660), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n664), .B1(new_n809), .B2(KEYINPUT102), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n658), .A2(new_n659), .A3(new_n660), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n671), .B1(new_n674), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n806), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n665), .A2(new_n672), .ZN(new_n817));
  OAI211_X1 g616(.A(KEYINPUT55), .B(new_n814), .C1(new_n665), .C2(new_n808), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n262), .A2(new_n245), .A3(new_n260), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n242), .B1(new_n241), .B2(new_n244), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n252), .A2(new_n253), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n259), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n820), .A2(new_n636), .A3(new_n642), .A4(new_n823), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n820), .B(new_n823), .C1(new_n673), .C2(new_n676), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n826), .B1(new_n819), .B2(new_n267), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n825), .B1(new_n827), .B2(new_n643), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n805), .B1(new_n828), .B2(new_n604), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT114), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n831), .B(new_n805), .C1(new_n828), .C2(new_n604), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n696), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n834), .A2(new_n683), .A3(new_n557), .A4(new_n556), .ZN(new_n835));
  OAI21_X1  g634(.A(G113gat), .B1(new_n835), .B2(new_n269), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n833), .A2(new_n682), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n536), .A2(new_n537), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n839), .A2(new_n686), .A3(new_n696), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n264), .A2(new_n271), .A3(new_n273), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n836), .B1(new_n841), .B2(new_n842), .ZN(G1340gat));
  NOR3_X1   g642(.A1(new_n835), .A2(new_n309), .A3(new_n677), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n837), .A2(new_n678), .A3(new_n840), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n309), .B2(new_n845), .ZN(G1341gat));
  OAI21_X1  g645(.A(G127gat), .B1(new_n835), .B2(new_n701), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n701), .A2(G127gat), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n841), .B2(new_n848), .ZN(G1342gat));
  NOR4_X1   g648(.A1(new_n841), .A2(new_n304), .A3(new_n305), .A4(new_n643), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n850), .B(KEYINPUT56), .ZN(new_n851));
  OAI21_X1  g650(.A(G134gat), .B1(new_n835), .B2(new_n643), .ZN(new_n852));
  XNOR2_X1  g651(.A(new_n852), .B(KEYINPUT115), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(G1343gat));
  NOR3_X1   g653(.A1(new_n736), .A2(new_n682), .A3(new_n686), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n498), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  AND2_X1   g658(.A1(new_n816), .A2(new_n817), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n266), .A2(new_n268), .A3(new_n818), .A4(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n715), .B1(new_n861), .B2(new_n826), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n701), .B1(new_n862), .B2(new_n825), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n859), .B1(new_n863), .B2(new_n805), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n830), .A2(new_n696), .A3(new_n832), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n857), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n864), .B1(new_n866), .B2(KEYINPUT116), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT116), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n865), .A2(new_n868), .A3(new_n857), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n856), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n286), .B1(new_n870), .B2(new_n264), .ZN(new_n871));
  INV_X1    g670(.A(new_n837), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n543), .A2(new_n696), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT117), .Z(new_n874));
  NOR2_X1   g673(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n686), .A2(new_n269), .A3(G141gat), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n871), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT58), .ZN(new_n878));
  INV_X1    g677(.A(new_n269), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n286), .B1(new_n870), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n875), .A2(KEYINPUT118), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n269), .A2(G141gat), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n883), .B1(new_n872), .B2(new_n874), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n881), .A2(new_n556), .A3(new_n882), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n878), .ZN(new_n886));
  OAI22_X1  g685(.A1(new_n877), .A2(new_n878), .B1(new_n880), .B2(new_n886), .ZN(G1344gat));
  XNOR2_X1  g686(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n679), .A2(new_n269), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n863), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT57), .B1(new_n890), .B2(new_n696), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n833), .A2(new_n859), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g692(.A1(new_n893), .A2(new_n678), .A3(new_n855), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n888), .B1(new_n894), .B2(new_n288), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n866), .A2(KEYINPUT116), .ZN(new_n896));
  INV_X1    g695(.A(new_n864), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n896), .A2(new_n869), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n678), .A3(new_n855), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n288), .A2(KEYINPUT59), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n899), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n895), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n881), .A2(new_n556), .A3(new_n884), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n905), .A2(new_n288), .A3(new_n678), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n904), .A2(new_n906), .ZN(G1345gat));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n291), .A3(new_n604), .ZN(new_n908));
  INV_X1    g707(.A(new_n870), .ZN(new_n909));
  OAI21_X1  g708(.A(G155gat), .B1(new_n909), .B2(new_n701), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n908), .A2(new_n910), .ZN(G1346gat));
  NOR3_X1   g710(.A1(new_n909), .A2(new_n292), .A3(new_n643), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n905), .A2(new_n715), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(new_n292), .ZN(G1347gat));
  NAND3_X1  g713(.A1(new_n834), .A2(new_n682), .A3(new_n686), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n915), .A2(new_n839), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n361), .A3(new_n264), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n915), .A2(new_n693), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n361), .B1(new_n918), .B2(new_n879), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT121), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n919), .A2(new_n920), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n917), .B1(new_n921), .B2(new_n922), .ZN(G1348gat));
  INV_X1    g722(.A(new_n918), .ZN(new_n924));
  OAI21_X1  g723(.A(G176gat), .B1(new_n924), .B2(new_n677), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n916), .A2(new_n362), .A3(new_n678), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(G1349gat));
  OAI21_X1  g726(.A(G183gat), .B1(new_n924), .B2(new_n701), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n701), .A2(new_n410), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n916), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g730(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n928), .A2(new_n930), .A3(new_n932), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1350gat));
  NAND3_X1  g735(.A1(new_n916), .A2(new_n379), .A3(new_n715), .ZN(new_n937));
  NAND2_X1  g736(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G190gat), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n939), .B1(new_n918), .B2(new_n715), .ZN(new_n940));
  NOR2_X1   g739(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n940), .A2(new_n941), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n937), .B1(new_n942), .B2(new_n943), .ZN(G1351gat));
  NOR3_X1   g743(.A1(new_n736), .A2(new_n683), .A3(new_n556), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n893), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(G197gat), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n946), .A2(new_n947), .A3(new_n269), .ZN(new_n948));
  INV_X1    g747(.A(new_n865), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n264), .A3(new_n945), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n948), .B1(new_n947), .B2(new_n950), .ZN(G1352gat));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n945), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n952), .A2(G204gat), .A3(new_n677), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT124), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n953), .A2(new_n954), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(G204gat), .B1(new_n946), .B2(new_n677), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n955), .A2(KEYINPUT62), .A3(new_n956), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(G1353gat));
  NAND4_X1  g761(.A1(new_n949), .A2(new_n432), .A3(new_n604), .A4(new_n945), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n945), .B(new_n604), .C1(new_n891), .C2(new_n892), .ZN(new_n964));
  AND3_X1   g763(.A1(new_n964), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n965));
  AOI21_X1  g764(.A(KEYINPUT63), .B1(new_n964), .B2(G211gat), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n963), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n967), .A2(KEYINPUT125), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n969));
  OAI211_X1 g768(.A(new_n969), .B(new_n963), .C1(new_n965), .C2(new_n966), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n968), .A2(new_n970), .ZN(G1354gat));
  OAI21_X1  g770(.A(new_n428), .B1(new_n952), .B2(new_n643), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT126), .Z(new_n973));
  INV_X1    g772(.A(new_n946), .ZN(new_n974));
  AOI211_X1 g773(.A(new_n431), .B(new_n643), .C1(new_n974), .C2(KEYINPUT127), .ZN(new_n975));
  OR2_X1    g774(.A1(new_n974), .A2(KEYINPUT127), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G1355gat));
endmodule


