//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:32 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n456, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n551, new_n552,
    new_n553, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  AOI22_X1  g029(.A1(new_n451), .A2(G2106), .B1(G567), .B2(new_n452), .ZN(G319));
  INV_X1    g030(.A(G2105), .ZN(new_n456));
  INV_X1    g031(.A(G137), .ZN(new_n457));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n458));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n457), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND2_X1   g037(.A1(G101), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n456), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n465), .B1(new_n460), .B2(new_n461), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(KEYINPUT65), .A2(G113), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G2105), .B1(new_n466), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n464), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n456), .ZN(new_n476));
  XNOR2_X1  g051(.A(new_n476), .B(KEYINPUT66), .ZN(new_n477));
  AND2_X1   g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NOR2_X1   g053(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n456), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(G2105), .ZN(new_n482));
  AOI22_X1  g057(.A1(G124), .A2(new_n481), .B1(new_n482), .B2(G136), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n477), .A2(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G138), .B(new_n456), .C1(new_n478), .C2(new_n479), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(KEYINPUT67), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT3), .B(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n491), .B1(new_n492), .B2(G126), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n489), .B1(new_n493), .B2(new_n456), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  AOI21_X1  g072(.A(new_n497), .B1(KEYINPUT67), .B2(new_n486), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n492), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(G102), .A2(G2104), .ZN(new_n500));
  AOI21_X1  g075(.A(G2105), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n494), .A2(new_n501), .ZN(G164));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(G50), .A3(G543), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT68), .ZN(new_n509));
  XNOR2_X1  g084(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  AOI21_X1  g086(.A(KEYINPUT69), .B1(KEYINPUT70), .B2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT69), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n504), .A2(new_n506), .ZN(new_n517));
  NOR3_X1   g092(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g093(.A(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n510), .B1(new_n511), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n515), .A2(new_n516), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n522), .A2(new_n503), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n520), .A2(new_n523), .ZN(G166));
  NAND2_X1  g099(.A1(new_n518), .A2(G89), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n526));
  AND3_X1   g101(.A1(new_n504), .A2(new_n506), .A3(G543), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n527), .A2(G51), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n525), .A2(new_n526), .A3(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(new_n521), .ZN(new_n535));
  INV_X1    g110(.A(G64), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n503), .B1(new_n537), .B2(KEYINPUT71), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n538), .B1(KEYINPUT71), .B2(new_n537), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n518), .A2(G90), .B1(G52), .B2(new_n527), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n518), .A2(G81), .B1(G43), .B2(new_n527), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT72), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n503), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT8), .ZN(new_n552));
  NAND4_X1  g127(.A1(G319), .A2(G483), .A3(G661), .A4(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT73), .ZN(G188));
  AND2_X1   g129(.A1(new_n513), .A2(new_n514), .ZN(new_n555));
  INV_X1    g130(.A(new_n516), .ZN(new_n556));
  AND3_X1   g131(.A1(new_n555), .A2(G65), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(G78), .A2(G543), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT74), .ZN(new_n562));
  INV_X1    g137(.A(new_n527), .ZN(new_n563));
  OAI21_X1  g138(.A(G53), .B1(new_n561), .B2(KEYINPUT74), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n527), .A2(KEYINPUT74), .A3(new_n561), .A4(G53), .ZN(new_n566));
  AOI22_X1  g141(.A1(new_n565), .A2(new_n566), .B1(new_n518), .B2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n560), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT75), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n568), .B(new_n569), .ZN(G299));
  INV_X1    g145(.A(G166), .ZN(G303));
  OAI21_X1  g146(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n521), .A2(G87), .A3(new_n507), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n527), .A2(G49), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  NAND3_X1  g150(.A1(new_n555), .A2(G61), .A3(new_n556), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n521), .A2(KEYINPUT76), .A3(G61), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n518), .A2(G86), .B1(G48), .B2(new_n527), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G305));
  AOI22_X1  g159(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n503), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n527), .A2(G47), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n519), .B2(new_n588), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(new_n518), .A2(G92), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT10), .Z(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n535), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n596), .A2(G651), .B1(G54), .B2(new_n527), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G171), .B2(new_n599), .ZN(G284));
  OAI21_X1  g176(.A(new_n600), .B1(G171), .B2(new_n599), .ZN(G321));
  NOR2_X1   g177(.A1(G286), .A2(new_n599), .ZN(new_n603));
  XNOR2_X1  g178(.A(G299), .B(KEYINPUT77), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(new_n599), .ZN(G297));
  AOI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(new_n599), .ZN(G280));
  AND2_X1   g181(.A1(new_n593), .A2(new_n597), .ZN(new_n607));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n548), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g188(.A1(new_n482), .A2(G2104), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  INV_X1    g191(.A(new_n616), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n617), .A2(G2100), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(KEYINPUT78), .Z(new_n619));
  NAND2_X1  g194(.A1(new_n482), .A2(G135), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n481), .A2(G123), .ZN(new_n621));
  NOR2_X1   g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(new_n456), .B2(G111), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2096), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n625), .B1(new_n617), .B2(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n619), .A2(new_n626), .ZN(G156));
  XNOR2_X1  g202(.A(G2451), .B(G2454), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT16), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT80), .ZN(new_n632));
  INV_X1    g207(.A(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G2427), .B(G2430), .Z(new_n635));
  NOR2_X1   g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT79), .B(KEYINPUT14), .ZN(new_n637));
  NOR2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT81), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n634), .A2(new_n635), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n639), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n641), .B1(new_n639), .B2(new_n642), .ZN(new_n645));
  OAI21_X1  g220(.A(new_n630), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  INV_X1    g221(.A(new_n645), .ZN(new_n647));
  NAND3_X1  g222(.A1(new_n647), .A2(new_n629), .A3(new_n643), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n646), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(KEYINPUT82), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g227(.A1(new_n646), .A2(new_n648), .A3(KEYINPUT82), .A4(new_n649), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g229(.A(new_n649), .B1(new_n646), .B2(new_n648), .ZN(new_n655));
  INV_X1    g230(.A(G14), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  XOR2_X1   g235(.A(G2084), .B(G2090), .Z(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(KEYINPUT83), .B(KEYINPUT18), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n660), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AND2_X1   g240(.A1(new_n663), .A2(KEYINPUT17), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n661), .A2(new_n662), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n664), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  MUX2_X1   g243(.A(new_n665), .B(new_n660), .S(new_n668), .Z(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT84), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n669), .B(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  NAND3_X1  g255(.A1(new_n675), .A2(new_n676), .A3(new_n677), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n676), .B(new_n677), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT85), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n680), .B(new_n681), .C1(new_n675), .C2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(G1991), .B(G1996), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT86), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1981), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n687), .B(new_n690), .ZN(G229));
  NAND2_X1  g266(.A1(KEYINPUT24), .A2(G34), .ZN(new_n692));
  INV_X1    g267(.A(KEYINPUT24), .ZN(new_n693));
  INV_X1    g268(.A(G34), .ZN(new_n694));
  AOI21_X1  g269(.A(G29), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI22_X1  g270(.A1(new_n473), .A2(G29), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G2084), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT96), .ZN(new_n699));
  AOI22_X1  g274(.A1(G129), .A2(new_n481), .B1(new_n482), .B2(G141), .ZN(new_n700));
  NAND3_X1  g275(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT26), .Z(new_n702));
  NAND3_X1  g277(.A1(new_n456), .A2(G105), .A3(G2104), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  MUX2_X1   g279(.A(G32), .B(new_n704), .S(G29), .Z(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT27), .B(G1996), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n708), .A2(G33), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT25), .ZN(new_n710));
  NAND2_X1  g285(.A1(G103), .A2(G2104), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(G2105), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n456), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n482), .A2(G139), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n456), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n709), .B1(new_n716), .B2(G29), .ZN(new_n717));
  XNOR2_X1  g292(.A(KEYINPUT94), .B(G2072), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n696), .A2(new_n697), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n482), .A2(G140), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n481), .A2(G128), .ZN(new_n723));
  NOR2_X1   g298(.A1(G104), .A2(G2105), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(new_n456), .B2(G116), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n722), .B(new_n723), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G29), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n708), .A2(G26), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT93), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT28), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G2067), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G28), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(KEYINPUT30), .ZN(new_n735));
  AOI21_X1  g310(.A(G29), .B1(new_n734), .B2(KEYINPUT30), .ZN(new_n736));
  OR2_X1    g311(.A1(KEYINPUT31), .A2(G11), .ZN(new_n737));
  NAND2_X1  g312(.A1(KEYINPUT31), .A2(G11), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n735), .A2(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n624), .B2(new_n708), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(new_n717), .B2(new_n718), .ZN(new_n741));
  NAND4_X1  g316(.A1(new_n707), .A2(new_n721), .A3(new_n733), .A4(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G21), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G168), .B2(new_n743), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n699), .B(new_n742), .C1(G1966), .C2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n708), .A2(G27), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G164), .B2(new_n708), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT97), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(G2078), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n745), .A2(G1966), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT95), .Z(new_n752));
  NOR2_X1   g327(.A1(new_n607), .A2(new_n743), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G4), .B2(new_n743), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT92), .B(G1348), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AND4_X1   g331(.A1(new_n746), .A2(new_n750), .A3(new_n752), .A4(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G171), .A2(new_n743), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G5), .B2(new_n743), .ZN(new_n759));
  INV_X1    g334(.A(G1961), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n743), .A2(G19), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n548), .B2(new_n743), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(G1341), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n743), .A2(G20), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT23), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n568), .B(KEYINPUT75), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(new_n743), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(G1956), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n708), .A2(G35), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n772), .B1(G162), .B2(new_n708), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT98), .Z(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT29), .ZN(new_n775));
  INV_X1    g350(.A(G2090), .ZN(new_n776));
  AND2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n754), .A2(new_n755), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n777), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n757), .A2(new_n765), .A3(new_n771), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G16), .A2(G24), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n590), .B(KEYINPUT88), .ZN(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1986), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT89), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n784), .A2(new_n785), .ZN(new_n788));
  AND3_X1   g363(.A1(new_n786), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n787), .B1(new_n786), .B2(new_n788), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n481), .A2(G119), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT87), .Z(new_n792));
  OR2_X1    g367(.A1(G95), .A2(G2105), .ZN(new_n793));
  INV_X1    g368(.A(G107), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n459), .B1(new_n794), .B2(G2105), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n482), .A2(G131), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  MUX2_X1   g372(.A(G25), .B(new_n797), .S(G29), .Z(new_n798));
  XOR2_X1   g373(.A(KEYINPUT35), .B(G1991), .Z(new_n799));
  INV_X1    g374(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n798), .B(new_n800), .ZN(new_n801));
  NOR3_X1   g376(.A1(new_n789), .A2(new_n790), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n743), .A2(G22), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G166), .B2(new_n743), .ZN(new_n804));
  XOR2_X1   g379(.A(KEYINPUT91), .B(G1971), .Z(new_n805));
  XOR2_X1   g380(.A(new_n804), .B(new_n805), .Z(new_n806));
  MUX2_X1   g381(.A(G6), .B(G305), .S(G16), .Z(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT32), .B(G1981), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AND2_X1   g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NOR3_X1   g385(.A1(new_n806), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT90), .ZN(new_n812));
  NAND2_X1  g387(.A1(G288), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT90), .A4(new_n574), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  MUX2_X1   g390(.A(G23), .B(new_n815), .S(G16), .Z(new_n816));
  OR2_X1    g391(.A1(new_n816), .A2(KEYINPUT33), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(KEYINPUT33), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(G1976), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n817), .A2(G1976), .A3(new_n818), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n811), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n823), .A2(KEYINPUT34), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT34), .ZN(new_n825));
  NAND4_X1  g400(.A1(new_n811), .A2(new_n825), .A3(new_n821), .A4(new_n822), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n802), .A2(new_n824), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT36), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT36), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n802), .A2(new_n824), .A3(new_n829), .A4(new_n826), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n781), .B1(new_n828), .B2(new_n830), .ZN(G311));
  INV_X1    g406(.A(KEYINPUT99), .ZN(new_n832));
  XNOR2_X1  g407(.A(G311), .B(new_n832), .ZN(G150));
  NAND2_X1  g408(.A1(new_n518), .A2(G93), .ZN(new_n834));
  XOR2_X1   g409(.A(KEYINPUT100), .B(G55), .Z(new_n835));
  AOI22_X1  g410(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n836));
  OAI221_X1 g411(.A(new_n834), .B1(new_n563), .B2(new_n835), .C1(new_n836), .C2(new_n503), .ZN(new_n837));
  OR2_X1    g412(.A1(new_n547), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n547), .A2(new_n837), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT38), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n607), .A2(G559), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n841), .B(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT39), .ZN(new_n844));
  AOI21_X1  g419(.A(G860), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n844), .B2(new_n843), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n837), .A2(G860), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT37), .Z(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(G145));
  XNOR2_X1  g424(.A(new_n704), .B(new_n716), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(new_n726), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT101), .B1(new_n494), .B2(new_n501), .ZN(new_n852));
  OAI21_X1  g427(.A(G126), .B1(new_n478), .B2(new_n479), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n853), .A2(new_n490), .ZN(new_n854));
  AOI22_X1  g429(.A1(new_n854), .A2(G2105), .B1(new_n488), .B2(new_n485), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n496), .A2(new_n487), .A3(G138), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n500), .B1(new_n856), .B2(new_n480), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n857), .A2(new_n456), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT101), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n852), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n851), .B(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n797), .B(new_n615), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n482), .A2(G142), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n481), .A2(G130), .ZN(new_n865));
  NOR2_X1   g440(.A1(G106), .A2(G2105), .ZN(new_n866));
  OAI21_X1  g441(.A(G2104), .B1(new_n456), .B2(G118), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n864), .B(new_n865), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n863), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n862), .B(new_n869), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n624), .B(G160), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(G162), .ZN(new_n872));
  AOI21_X1  g447(.A(G37), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n862), .A2(new_n869), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(KEYINPUT102), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(KEYINPUT102), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n862), .A2(new_n869), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n877), .A2(new_n872), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT40), .Z(G395));
  XOR2_X1   g456(.A(new_n840), .B(new_n610), .Z(new_n882));
  NAND2_X1  g457(.A1(G299), .A2(new_n607), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n768), .A2(new_n598), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT41), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT41), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n882), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n885), .A2(KEYINPUT103), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n887), .A2(new_n893), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n891), .B1(new_n895), .B2(new_n882), .ZN(new_n896));
  OR2_X1    g471(.A1(new_n896), .A2(KEYINPUT42), .ZN(new_n897));
  XNOR2_X1  g472(.A(new_n815), .B(new_n590), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n898), .A2(KEYINPUT104), .ZN(new_n899));
  XOR2_X1   g474(.A(G305), .B(G166), .Z(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n898), .A2(KEYINPUT104), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(KEYINPUT104), .A3(new_n898), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n896), .A2(KEYINPUT42), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n897), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n905), .B1(new_n897), .B2(new_n906), .ZN(new_n908));
  OAI21_X1  g483(.A(G868), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n837), .A2(new_n599), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(G295));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n910), .ZN(G331));
  XNOR2_X1  g487(.A(G301), .B(G168), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(new_n840), .ZN(new_n914));
  INV_X1    g489(.A(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n840), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n890), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n916), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n887), .B1(new_n918), .B2(new_n914), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n905), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(G37), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n905), .B1(new_n917), .B2(new_n919), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT43), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n894), .B(new_n892), .C1(new_n918), .C2(new_n914), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n903), .A2(new_n904), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n889), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n915), .A2(new_n916), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n927), .B1(new_n886), .B2(new_n889), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n925), .B(new_n926), .C1(new_n929), .C2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n931), .A2(new_n920), .A3(new_n932), .A4(new_n921), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n924), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n934), .A2(KEYINPUT44), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n931), .A2(new_n920), .A3(new_n921), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(KEYINPUT43), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n940));
  OR3_X1    g515(.A1(new_n922), .A2(KEYINPUT43), .A3(new_n923), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n935), .B1(new_n942), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g518(.A(KEYINPUT125), .ZN(new_n944));
  XNOR2_X1  g519(.A(new_n726), .B(new_n732), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n704), .B(G1996), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n797), .A2(new_n800), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n797), .A2(new_n800), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(G290), .A2(G1986), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n590), .A2(new_n785), .ZN(new_n954));
  NOR3_X1   g529(.A1(new_n952), .A2(new_n953), .A3(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT45), .B1(new_n861), .B2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n464), .A2(new_n472), .A3(G40), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT107), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n464), .A2(new_n472), .A3(new_n960), .A4(G40), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n957), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n955), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n956), .B1(new_n494), .B2(new_n501), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(G1384), .ZN(new_n968));
  INV_X1    g543(.A(new_n968), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n967), .B(new_n962), .C1(G164), .C2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n971));
  OR3_X1    g546(.A1(new_n970), .A2(new_n971), .A3(G2078), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n852), .A2(new_n860), .A3(new_n968), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(new_n962), .A3(new_n967), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n971), .B1(new_n974), .B2(G2078), .ZN(new_n975));
  AOI21_X1  g550(.A(G1384), .B1(new_n855), .B2(new_n858), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT50), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n965), .A2(KEYINPUT50), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(new_n979), .A3(new_n962), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n760), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n972), .A2(new_n975), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(G171), .ZN(new_n983));
  AND2_X1   g558(.A1(new_n975), .A2(new_n981), .ZN(new_n984));
  NOR3_X1   g559(.A1(new_n958), .A2(new_n971), .A3(G2078), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n973), .A2(new_n985), .ZN(new_n986));
  OR3_X1    g561(.A1(new_n957), .A2(KEYINPUT123), .A3(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(KEYINPUT123), .B1(new_n957), .B2(new_n986), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n984), .A2(G301), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n983), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n984), .A2(G301), .A3(new_n972), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n984), .A2(new_n988), .A3(new_n987), .ZN(new_n994));
  OAI211_X1 g569(.A(KEYINPUT54), .B(new_n993), .C1(new_n994), .C2(G301), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT51), .ZN(new_n996));
  INV_X1    g571(.A(G8), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1966), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n970), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n980), .A2(G2084), .ZN(new_n1002));
  OAI21_X1  g577(.A(G168), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AND3_X1   g578(.A1(new_n978), .A2(new_n979), .A3(new_n962), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n697), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n970), .A2(new_n1000), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(G286), .A3(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n999), .B1(new_n1003), .B2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1005), .A2(G168), .A3(new_n1006), .ZN(new_n1009));
  AOI21_X1  g584(.A(KEYINPUT51), .B1(new_n1009), .B2(G8), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n992), .A2(new_n995), .A3(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(KEYINPUT108), .B(G2090), .ZN(new_n1013));
  INV_X1    g588(.A(G1971), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1004), .A2(new_n1013), .B1(new_n974), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT109), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT109), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n974), .A2(new_n1014), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1013), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n980), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1017), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(G8), .B1(new_n520), .B2(new_n523), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT55), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1022), .B(new_n1023), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1016), .A2(new_n1021), .A3(G8), .A4(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(new_n1022), .B(KEYINPUT55), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1026), .B1(new_n997), .B2(new_n1015), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(G288), .A2(new_n820), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1030), .A2(KEYINPUT52), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n965), .B1(new_n961), .B2(new_n959), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n1032), .A2(new_n997), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n813), .A2(G1976), .A3(new_n814), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1036), .B1(new_n1037), .B2(KEYINPUT52), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n1039));
  AOI211_X1 g614(.A(KEYINPUT110), .B(new_n1039), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1035), .B1(new_n1038), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT112), .ZN(new_n1042));
  INV_X1    g617(.A(G1981), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n582), .A2(new_n1043), .A3(new_n583), .ZN(new_n1044));
  INV_X1    g619(.A(new_n580), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n576), .B2(new_n577), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n503), .B1(new_n1046), .B2(new_n579), .ZN(new_n1047));
  INV_X1    g622(.A(new_n583), .ZN(new_n1048));
  OAI21_X1  g623(.A(G1981), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT49), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(KEYINPUT111), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1044), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n1033), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1051), .B1(new_n1044), .B2(new_n1049), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1042), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1044), .A2(new_n1049), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1056), .A2(KEYINPUT111), .A3(new_n1050), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n1057), .A2(KEYINPUT112), .A3(new_n1033), .A4(new_n1052), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1041), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT124), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1029), .A2(new_n1059), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1055), .A2(new_n1058), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1035), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1037), .A2(KEYINPUT52), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(KEYINPUT110), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1037), .A2(new_n1036), .A3(KEYINPUT52), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1063), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1062), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(KEYINPUT124), .B1(new_n1068), .B2(new_n1028), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1012), .B1(new_n1061), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT60), .ZN(new_n1071));
  INV_X1    g646(.A(new_n755), .ZN(new_n1072));
  AOI22_X1  g647(.A1(KEYINPUT50), .A2(new_n965), .B1(new_n959), .B2(new_n961), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1072), .B1(new_n1073), .B2(new_n978), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n962), .A2(new_n732), .A3(new_n976), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT116), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT116), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1078), .B(new_n1075), .C1(new_n1004), .C2(new_n1072), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1071), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1077), .A2(new_n1071), .A3(new_n1079), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1082), .A2(new_n1083), .A3(new_n607), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1083), .B1(new_n1082), .B2(new_n607), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1081), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1082), .A2(new_n607), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(KEYINPUT122), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1082), .A2(new_n1083), .A3(new_n607), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1088), .A2(new_n1080), .A3(new_n1089), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1092), .B1(new_n560), .B2(new_n567), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n560), .A2(new_n567), .A3(new_n1092), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(G1956), .B1(new_n1073), .B2(new_n978), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT56), .B(G2072), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n962), .A2(new_n973), .A3(new_n967), .A4(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1096), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1956), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n980), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n973), .A2(new_n967), .A3(new_n962), .A4(new_n1098), .ZN(new_n1103));
  NAND4_X1  g678(.A1(new_n1102), .A2(new_n1094), .A3(new_n1095), .A4(new_n1103), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1100), .A2(KEYINPUT61), .A3(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT120), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1100), .A2(new_n1104), .A3(KEYINPUT120), .A4(KEYINPUT61), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT119), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT58), .B(G1341), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1110), .B1(new_n1032), .B2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n962), .A2(new_n976), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1111), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1113), .A2(KEYINPUT119), .A3(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g690(.A(KEYINPUT118), .B(G1996), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n973), .A2(new_n967), .A3(new_n962), .A4(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1112), .A2(new_n1115), .A3(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n548), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(KEYINPUT59), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT59), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1118), .A2(new_n548), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT61), .ZN(new_n1124));
  AOI22_X1  g699(.A1(new_n1120), .A2(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  AND3_X1   g700(.A1(new_n1109), .A2(KEYINPUT121), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(KEYINPUT121), .B1(new_n1109), .B2(new_n1125), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1091), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1077), .A2(new_n607), .A3(new_n1079), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT117), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1100), .B1(new_n1129), .B2(KEYINPUT117), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(new_n1104), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1070), .B1(new_n1128), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(new_n1033), .ZN(new_n1137));
  NOR2_X1   g712(.A1(G288), .A2(G1976), .ZN(new_n1138));
  XNOR2_X1  g713(.A(new_n1138), .B(KEYINPUT114), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1062), .A2(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n1044), .B(KEYINPUT113), .Z(new_n1141));
  AOI21_X1  g716(.A(new_n1137), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(G286), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1144), .A2(KEYINPUT63), .A3(G8), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1016), .A2(new_n1021), .A3(G8), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1026), .ZN(new_n1147));
  AND4_X1   g722(.A1(new_n1059), .A2(new_n1025), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT115), .B(KEYINPUT63), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n974), .A2(new_n1014), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1150), .B1(new_n980), .B2(new_n1019), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1144), .B(G8), .C1(new_n1024), .C2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1025), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1149), .B1(new_n1059), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1143), .B1(new_n1148), .B2(new_n1154), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1005), .A2(G286), .A3(new_n1006), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n998), .B1(new_n1156), .B2(new_n1144), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1009), .A2(G8), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1157), .B(KEYINPUT62), .C1(KEYINPUT51), .C2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1160), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1161));
  INV_X1    g736(.A(new_n983), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1163), .B1(new_n1061), .B2(new_n1069), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1155), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n964), .B1(new_n1136), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g741(.A1(new_n963), .A2(G1996), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n1167), .A2(KEYINPUT46), .ZN(new_n1168));
  INV_X1    g743(.A(new_n963), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1169), .B1(new_n704), .B2(new_n946), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1171), .B1(KEYINPUT46), .B2(new_n1167), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1172), .A2(KEYINPUT47), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1172), .A2(KEYINPUT47), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT48), .B1(new_n1169), .B2(new_n953), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1175), .B1(new_n1169), .B2(new_n952), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1169), .A2(KEYINPUT48), .A3(new_n953), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n948), .A2(new_n949), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(G2067), .B2(new_n726), .ZN(new_n1179));
  AOI22_X1  g754(.A1(new_n1176), .A2(new_n1177), .B1(new_n1169), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1173), .A2(new_n1174), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n944), .B1(new_n1166), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1181), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1060), .B1(new_n1029), .B2(new_n1059), .ZN(new_n1185));
  NOR3_X1   g760(.A1(new_n1068), .A2(new_n1028), .A3(KEYINPUT124), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(new_n1149), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1153), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1188), .B1(new_n1189), .B2(new_n1068), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1059), .A2(new_n1145), .A3(new_n1025), .A4(new_n1147), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1142), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1187), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1127), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1109), .A2(new_n1125), .A3(KEYINPUT121), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1134), .B1(new_n1196), .B2(new_n1091), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1193), .B1(new_n1197), .B2(new_n1070), .ZN(new_n1198));
  OAI211_X1 g773(.A(KEYINPUT125), .B(new_n1183), .C1(new_n1198), .C2(new_n964), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1182), .A2(new_n1199), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g775(.A1(new_n880), .A2(G229), .ZN(new_n1202));
  NAND2_X1  g776(.A1(new_n672), .A2(G319), .ZN(new_n1203));
  XNOR2_X1  g777(.A(new_n1203), .B(KEYINPUT126), .ZN(new_n1204));
  INV_X1    g778(.A(new_n1204), .ZN(new_n1205));
  AOI21_X1  g779(.A(KEYINPUT127), .B1(new_n658), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n1207));
  AOI211_X1 g781(.A(new_n1207), .B(new_n1204), .C1(new_n654), .C2(new_n657), .ZN(new_n1208));
  OAI211_X1 g782(.A(new_n934), .B(new_n1202), .C1(new_n1206), .C2(new_n1208), .ZN(G225));
  INV_X1    g783(.A(G225), .ZN(G308));
endmodule


