//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:35 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n744, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1069, new_n1070, new_n1071, new_n1072,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT9), .B(G234), .Z(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n188), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(G110), .B(G140), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  AND2_X1   g007(.A1(new_n193), .A2(G227), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n192), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT78), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT10), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT76), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G146), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(new_n203), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(KEYINPUT67), .ZN(new_n207));
  XNOR2_X1  g021(.A(G143), .B(G146), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(new_n201), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n207), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g025(.A(KEYINPUT1), .B1(new_n204), .B2(G146), .ZN(new_n212));
  AOI22_X1  g026(.A1(new_n212), .A2(G128), .B1(new_n203), .B2(new_n205), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G104), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT3), .B1(new_n216), .B2(G107), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G104), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(G107), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n217), .A2(new_n220), .A3(new_n221), .A4(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n216), .A2(G107), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n219), .A2(G104), .ZN(new_n225));
  OAI21_X1  g039(.A(G101), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n199), .B1(new_n215), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n213), .B1(new_n207), .B2(new_n210), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n230), .A2(KEYINPUT76), .A3(new_n227), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n198), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n204), .A2(KEYINPUT64), .A3(G146), .ZN(new_n233));
  AOI21_X1  g047(.A(KEYINPUT64), .B1(new_n204), .B2(G146), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n203), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n212), .A2(G128), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n235), .A2(KEYINPUT68), .A3(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n204), .A2(G146), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT64), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n240), .B1(new_n202), .B2(G143), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n204), .A2(KEYINPUT64), .A3(G146), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n239), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n200), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n238), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n237), .A2(new_n245), .A3(new_n211), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n245), .A2(new_n237), .A3(new_n211), .A4(KEYINPUT70), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n227), .A2(new_n198), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n217), .A2(new_n220), .A3(new_n222), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G101), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n253), .A2(KEYINPUT4), .A3(new_n223), .ZN(new_n254));
  AND2_X1   g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  NOR2_X1   g069(.A1(KEYINPUT0), .A2(G128), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n235), .A2(new_n257), .B1(new_n208), .B2(new_n255), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n252), .A2(new_n259), .A3(G101), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n254), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n232), .A2(new_n251), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT77), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT11), .ZN(new_n265));
  INV_X1    g079(.A(G134), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(G137), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(G137), .ZN(new_n268));
  INV_X1    g082(.A(G137), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT11), .A3(G134), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G131), .ZN(new_n272));
  XNOR2_X1  g086(.A(KEYINPUT65), .B(G131), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n273), .A2(new_n267), .A3(new_n268), .A4(new_n270), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n232), .A2(new_n251), .A3(KEYINPUT77), .A4(new_n261), .ZN(new_n276));
  AND4_X1   g090(.A1(new_n197), .A2(new_n264), .A3(new_n275), .A4(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(new_n272), .A2(new_n274), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n232), .A2(new_n251), .A3(new_n278), .A4(new_n261), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT78), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n278), .B1(new_n262), .B2(new_n263), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n280), .B1(new_n281), .B2(new_n276), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n196), .B1(new_n277), .B2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n215), .A2(new_n199), .A3(new_n228), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT76), .B1(new_n230), .B2(new_n227), .ZN(new_n285));
  INV_X1    g099(.A(new_n246), .ZN(new_n286));
  AOI22_X1  g100(.A1(new_n284), .A2(new_n285), .B1(new_n286), .B2(new_n227), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT12), .B1(new_n287), .B2(new_n278), .ZN(new_n288));
  OAI22_X1  g102(.A1(new_n229), .A2(new_n231), .B1(new_n246), .B2(new_n228), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT12), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n289), .A2(new_n290), .A3(new_n275), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n288), .A2(new_n279), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n195), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n283), .A2(G469), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(G469), .A2(G902), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n264), .A2(new_n275), .A3(new_n276), .ZN(new_n297));
  INV_X1    g111(.A(new_n280), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n281), .A2(new_n197), .A3(new_n276), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n299), .A2(new_n195), .A3(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n292), .A2(new_n195), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI211_X1 g117(.A(G469), .B(G902), .C1(new_n301), .C2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n191), .B1(new_n296), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(G214), .B1(G237), .B2(G902), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  XOR2_X1   g121(.A(KEYINPUT2), .B(G113), .Z(new_n308));
  XNOR2_X1  g122(.A(G116), .B(G119), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G119), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G116), .ZN(new_n312));
  INV_X1    g126(.A(G116), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G119), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT2), .B(G113), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n310), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n254), .A2(new_n260), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G113), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n313), .A2(G119), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n320), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT5), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT79), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT5), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(new_n309), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n228), .A2(new_n310), .A3(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(KEYINPUT80), .B1(new_n319), .B2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n319), .A2(KEYINPUT80), .A3(new_n331), .ZN(new_n334));
  XNOR2_X1  g148(.A(G110), .B(G122), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n333), .A2(KEYINPUT6), .A3(new_n334), .A4(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT6), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n319), .A2(new_n331), .A3(new_n335), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT81), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n319), .A2(new_n331), .A3(KEYINPUT81), .A4(new_n335), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n338), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  AND3_X1   g157(.A1(new_n319), .A2(KEYINPUT80), .A3(new_n331), .ZN(new_n344));
  NOR3_X1   g158(.A1(new_n344), .A2(new_n332), .A3(new_n335), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n337), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT82), .ZN(new_n347));
  INV_X1    g161(.A(G125), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n347), .B1(new_n258), .B2(new_n348), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n245), .A2(new_n237), .A3(new_n211), .A4(new_n348), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n208), .A2(new_n255), .ZN(new_n351));
  INV_X1    g165(.A(new_n257), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n351), .B1(new_n243), .B2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(KEYINPUT82), .A3(G125), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n349), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n193), .A2(G224), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n349), .A2(new_n350), .A3(new_n356), .A4(new_n354), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n346), .A2(new_n360), .ZN(new_n361));
  XOR2_X1   g175(.A(KEYINPUT84), .B(KEYINPUT7), .Z(new_n362));
  OAI21_X1  g176(.A(new_n355), .B1(new_n357), .B2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT85), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n355), .B(KEYINPUT85), .C1(new_n357), .C2(new_n362), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT7), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n359), .A2(new_n368), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n323), .A2(new_n329), .B1(new_n309), .B2(new_n308), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n310), .A2(new_n223), .A3(new_n226), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n322), .A2(new_n325), .A3(new_n327), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n312), .A2(new_n314), .A3(KEYINPUT5), .ZN(new_n373));
  AND3_X1   g187(.A1(new_n372), .A2(new_n373), .A3(G113), .ZN(new_n374));
  OAI22_X1  g188(.A1(new_n370), .A2(new_n228), .B1(new_n371), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT83), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n335), .B(KEYINPUT8), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n376), .B1(new_n375), .B2(new_n377), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n369), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n341), .A2(new_n342), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n367), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n361), .A2(new_n189), .A3(new_n382), .ZN(new_n383));
  OAI21_X1  g197(.A(G210), .B1(G237), .B2(G902), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(KEYINPUT86), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(new_n385), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n361), .A2(new_n382), .A3(new_n189), .A4(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n307), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n305), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT32), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT31), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n269), .A2(G134), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(new_n268), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G131), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n274), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n248), .A2(new_n249), .A3(new_n397), .ZN(new_n398));
  AND3_X1   g212(.A1(new_n258), .A2(KEYINPUT69), .A3(new_n275), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT69), .B1(new_n258), .B2(new_n275), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n398), .A2(KEYINPUT30), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n246), .A2(new_n397), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT66), .B1(new_n278), .B2(new_n353), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT66), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n258), .A2(new_n275), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT30), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n402), .A2(new_n318), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n318), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n398), .A2(new_n411), .A3(new_n401), .ZN(new_n412));
  NOR2_X1   g226(.A1(G237), .A2(G953), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G210), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT27), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT26), .B(G101), .ZN(new_n416));
  XNOR2_X1  g230(.A(new_n415), .B(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n412), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n393), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n412), .A2(new_n417), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n402), .A2(new_n318), .A3(new_n409), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(KEYINPUT31), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n407), .A2(new_n318), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n412), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT28), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n318), .B1(new_n258), .B2(new_n275), .ZN(new_n426));
  AOI21_X1  g240(.A(KEYINPUT28), .B1(new_n398), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(new_n417), .ZN(new_n430));
  AOI22_X1  g244(.A1(new_n419), .A2(new_n422), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(G472), .A2(G902), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n392), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT28), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(new_n412), .B2(new_n423), .ZN(new_n436));
  NOR3_X1   g250(.A1(new_n436), .A2(new_n427), .A3(new_n430), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n417), .B1(new_n421), .B2(new_n412), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n437), .A2(new_n438), .A3(KEYINPUT29), .ZN(new_n439));
  INV_X1    g253(.A(new_n412), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n411), .B1(new_n398), .B2(new_n401), .ZN(new_n441));
  OAI21_X1  g255(.A(KEYINPUT28), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT29), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n430), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(new_n428), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n189), .ZN(new_n446));
  OAI21_X1  g260(.A(G472), .B1(new_n439), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n430), .B1(new_n436), .B2(new_n427), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n420), .A2(KEYINPUT31), .A3(new_n421), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT31), .B1(new_n420), .B2(new_n421), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n448), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT32), .A3(new_n432), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n434), .A2(new_n447), .A3(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT22), .B(G137), .ZN(new_n454));
  INV_X1    g268(.A(G234), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n187), .A2(new_n455), .A3(G953), .ZN(new_n456));
  XOR2_X1   g270(.A(new_n454), .B(new_n456), .Z(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G140), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G125), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n348), .A2(G140), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT16), .ZN(new_n462));
  OR3_X1    g276(.A1(new_n348), .A2(KEYINPUT16), .A3(G140), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n202), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(new_n463), .A3(G146), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n200), .A2(G119), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n311), .A2(G128), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT24), .B(G110), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT73), .ZN(new_n473));
  OAI21_X1  g287(.A(KEYINPUT23), .B1(new_n200), .B2(G119), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT71), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT71), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n469), .A2(new_n476), .A3(KEYINPUT23), .ZN(new_n477));
  OR3_X1    g291(.A1(new_n311), .A2(KEYINPUT72), .A3(G128), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n468), .A2(KEYINPUT72), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n475), .A2(new_n477), .A3(new_n478), .A4(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n200), .A2(KEYINPUT23), .A3(G119), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n473), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(G110), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n480), .A2(new_n473), .A3(new_n481), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n472), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n480), .A2(new_n483), .A3(new_n481), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n470), .A2(new_n471), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n460), .A2(new_n461), .A3(new_n202), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT74), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n460), .A2(new_n461), .A3(KEYINPUT74), .A4(new_n202), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n489), .A2(new_n466), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n458), .B1(new_n486), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n485), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n498), .A2(new_n482), .A3(new_n483), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n495), .B(new_n457), .C1(new_n499), .C2(new_n472), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(new_n500), .A3(new_n189), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT75), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT25), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(G217), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n505), .B1(G234), .B2(new_n189), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n501), .A2(new_n503), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n497), .A2(new_n500), .A3(KEYINPUT25), .A4(new_n189), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(KEYINPUT75), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n506), .A2(G902), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n497), .A2(new_n500), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(G475), .ZN(new_n516));
  INV_X1    g330(.A(G237), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n193), .A3(G214), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n204), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n413), .A2(G143), .A3(G214), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(KEYINPUT18), .A2(G131), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n521), .B(new_n522), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n202), .B1(new_n460), .B2(new_n461), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT87), .B1(new_n494), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT87), .ZN(new_n527));
  AOI211_X1 g341(.A(new_n527), .B(new_n524), .C1(new_n492), .C2(new_n493), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n523), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  XOR2_X1   g343(.A(KEYINPUT65), .B(G131), .Z(new_n530));
  OAI21_X1  g344(.A(KEYINPUT88), .B1(new_n521), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT17), .ZN(new_n532));
  INV_X1    g346(.A(new_n520), .ZN(new_n533));
  AOI21_X1  g347(.A(G143), .B1(new_n413), .B2(G214), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n530), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT88), .ZN(new_n536));
  NAND4_X1  g350(.A1(new_n519), .A2(new_n536), .A3(new_n273), .A4(new_n520), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n531), .A2(new_n532), .A3(new_n535), .A4(new_n537), .ZN(new_n538));
  OAI211_X1 g352(.A(KEYINPUT17), .B(new_n530), .C1(new_n533), .C2(new_n534), .ZN(new_n539));
  AND3_X1   g353(.A1(new_n539), .A2(new_n465), .A3(new_n466), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(G113), .B(G122), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(new_n216), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n529), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n543), .B1(new_n529), .B2(new_n541), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n189), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n516), .B1(new_n546), .B2(KEYINPUT90), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT90), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n548), .B(new_n189), .C1(new_n544), .C2(new_n545), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(G475), .A2(G902), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n533), .A2(new_n534), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n536), .B1(new_n552), .B2(new_n273), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n535), .A2(new_n537), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT89), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT89), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n531), .A2(new_n556), .A3(new_n535), .A4(new_n537), .ZN(new_n557));
  INV_X1    g371(.A(new_n466), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n460), .A2(new_n461), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT19), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n558), .B1(new_n561), .B2(new_n202), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n555), .A2(new_n557), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n543), .B1(new_n563), .B2(new_n529), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n551), .B1(new_n564), .B2(new_n544), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT20), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT20), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n567), .B(new_n551), .C1(new_n564), .C2(new_n544), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G478), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n570), .A2(KEYINPUT15), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT92), .ZN(new_n573));
  INV_X1    g387(.A(G122), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G116), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n313), .A2(G122), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n219), .ZN(new_n578));
  XNOR2_X1  g392(.A(G116), .B(G122), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(G107), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n204), .A2(G128), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n200), .A2(G143), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT13), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT13), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n204), .A3(G128), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G134), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n578), .B(new_n580), .C1(new_n583), .C2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n581), .A2(new_n582), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT91), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT91), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n581), .A2(new_n582), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(G134), .B1(new_n589), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n573), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n578), .A2(new_n580), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n581), .A2(new_n582), .A3(new_n590), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n590), .B1(new_n581), .B2(new_n582), .ZN(new_n596));
  OAI21_X1  g410(.A(new_n266), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(G134), .B(new_n585), .C1(new_n588), .C2(new_n584), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n594), .A2(new_n597), .A3(KEYINPUT92), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n589), .A2(G134), .A3(new_n591), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n219), .B1(new_n575), .B2(KEYINPUT14), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(new_n579), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n188), .A2(G217), .A3(new_n193), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n607), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n600), .A2(new_n605), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n572), .B1(new_n611), .B2(new_n189), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n600), .A2(new_n605), .A3(new_n609), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n609), .B1(new_n600), .B2(new_n605), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n189), .B(new_n572), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  OAI211_X1 g431(.A(G902), .B(G953), .C1(new_n455), .C2(new_n517), .ZN(new_n618));
  XOR2_X1   g432(.A(new_n618), .B(KEYINPUT94), .Z(new_n619));
  XNOR2_X1  g433(.A(KEYINPUT21), .B(G898), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(KEYINPUT93), .A2(G952), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(KEYINPUT93), .A2(G952), .ZN(new_n624));
  AOI21_X1  g438(.A(G953), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n625), .B1(new_n455), .B2(new_n517), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n550), .A2(new_n569), .A3(new_n617), .A4(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT95), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AOI22_X1  g444(.A1(new_n547), .A2(new_n549), .B1(new_n566), .B2(new_n568), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n631), .A2(KEYINPUT95), .A3(new_n627), .A4(new_n617), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n453), .A2(new_n515), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n391), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G101), .ZN(G3));
  NAND2_X1  g450(.A1(new_n451), .A2(new_n189), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n637), .A2(KEYINPUT96), .A3(G472), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n419), .A2(new_n422), .ZN(new_n639));
  AOI21_X1  g453(.A(G902), .B1(new_n639), .B2(new_n448), .ZN(new_n640));
  NAND2_X1  g454(.A1(KEYINPUT96), .A2(G472), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  NOR3_X1   g457(.A1(new_n305), .A2(new_n643), .A3(new_n514), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n306), .B1(new_n388), .B2(KEYINPUT97), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n386), .A2(KEYINPUT97), .A3(new_n388), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(new_n647), .A3(new_n627), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n613), .A2(new_n614), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(G902), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT100), .B(G478), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT99), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT33), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n654), .B1(new_n611), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n650), .A2(KEYINPUT99), .A3(KEYINPUT33), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n655), .B1(new_n613), .B2(new_n614), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(KEYINPUT98), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT98), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n611), .A2(new_n660), .A3(new_n655), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n656), .A2(new_n657), .B1(new_n659), .B2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n570), .A2(G902), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n653), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n649), .B1(new_n664), .B2(new_n631), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n656), .A2(new_n657), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n659), .A2(new_n661), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n666), .A2(new_n667), .A3(new_n663), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n668), .B1(new_n651), .B2(new_n652), .ZN(new_n669));
  INV_X1    g483(.A(new_n631), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(KEYINPUT101), .A3(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n648), .B1(new_n665), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n644), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT34), .B(G104), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G6));
  NOR2_X1   g489(.A1(new_n670), .A2(new_n617), .ZN(new_n676));
  AND4_X1   g490(.A1(new_n627), .A2(new_n646), .A3(new_n676), .A4(new_n647), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n644), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT102), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT35), .B(G107), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G9));
  NOR2_X1   g495(.A1(new_n486), .A2(new_n496), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n458), .A2(KEYINPUT36), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n684), .A2(new_n512), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n507), .B2(new_n510), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n630), .B2(new_n632), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n687), .A2(new_n642), .A3(new_n638), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n391), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT103), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT37), .B(G110), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G12));
  AND4_X1   g506(.A1(new_n189), .A2(new_n361), .A3(new_n387), .A4(new_n382), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n378), .A2(new_n379), .ZN(new_n694));
  AND2_X1   g508(.A1(new_n349), .A2(new_n354), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n695), .A2(KEYINPUT7), .A3(new_n356), .A4(new_n350), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n694), .A2(new_n381), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g511(.A(G902), .B1(new_n697), .B2(new_n367), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n387), .B1(new_n698), .B2(new_n361), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n693), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n645), .B1(new_n700), .B2(KEYINPUT97), .ZN(new_n701));
  INV_X1    g515(.A(new_n626), .ZN(new_n702));
  INV_X1    g516(.A(G900), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n702), .B1(new_n619), .B2(new_n703), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n670), .A2(new_n617), .A3(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n701), .A2(new_n453), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n684), .A2(new_n512), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n508), .A2(KEYINPUT75), .A3(new_n509), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n504), .A2(new_n506), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n707), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  OAI211_X1 g524(.A(new_n191), .B(new_n710), .C1(new_n296), .C2(new_n304), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n200), .ZN(G30));
  INV_X1    g527(.A(new_n293), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n299), .A2(new_n300), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n714), .B1(new_n715), .B2(new_n196), .ZN(new_n716));
  OAI21_X1  g530(.A(G469), .B1(new_n716), .B2(G902), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n301), .A2(new_n303), .ZN(new_n718));
  INV_X1    g532(.A(G469), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n718), .A2(new_n719), .A3(new_n189), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n190), .B1(new_n717), .B2(new_n720), .ZN(new_n721));
  XOR2_X1   g535(.A(new_n704), .B(KEYINPUT39), .Z(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n723), .A2(KEYINPUT40), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT104), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n398), .A2(new_n401), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n318), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(new_n412), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n189), .B1(new_n728), .B2(new_n417), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n430), .B1(new_n421), .B2(new_n412), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n725), .B(G472), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(G472), .B1(new_n729), .B2(new_n730), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(KEYINPUT104), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n434), .A2(new_n452), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT105), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n723), .A2(KEYINPUT40), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n386), .A2(new_n388), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT38), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n631), .A2(new_n617), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n306), .A3(new_n686), .A4(new_n740), .ZN(new_n741));
  NOR4_X1   g555(.A1(new_n724), .A2(new_n736), .A3(new_n737), .A4(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(new_n204), .ZN(G45));
  NOR3_X1   g557(.A1(new_n664), .A2(new_n631), .A3(new_n704), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n701), .A2(new_n453), .A3(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n711), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n202), .ZN(G48));
  AND2_X1   g561(.A1(new_n453), .A2(new_n515), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n719), .B1(new_n718), .B2(new_n189), .ZN(new_n749));
  NOR3_X1   g563(.A1(new_n749), .A2(new_n304), .A3(new_n190), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n665), .A2(new_n671), .ZN(new_n751));
  INV_X1    g565(.A(new_n648), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n748), .A2(new_n750), .A3(new_n751), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT41), .B(G113), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G15));
  NAND3_X1  g569(.A1(new_n748), .A2(new_n750), .A3(new_n677), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G116), .ZN(G18));
  INV_X1    g571(.A(KEYINPUT106), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n277), .A2(new_n282), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n302), .B1(new_n759), .B2(new_n195), .ZN(new_n760));
  OAI21_X1  g574(.A(G469), .B1(new_n760), .B2(G902), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n701), .A2(new_n191), .A3(new_n720), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n687), .A2(new_n453), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n758), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n687), .A2(new_n453), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(new_n750), .A3(KEYINPUT106), .A4(new_n701), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G119), .ZN(G21));
  INV_X1    g582(.A(KEYINPUT107), .ZN(new_n769));
  INV_X1    g583(.A(G472), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n769), .B1(new_n640), .B2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n637), .A2(KEYINPUT107), .A3(G472), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n427), .B1(new_n728), .B2(KEYINPUT28), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n639), .B1(new_n417), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n432), .ZN(new_n775));
  AND4_X1   g589(.A1(new_n515), .A2(new_n771), .A3(new_n772), .A4(new_n775), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n740), .A2(new_n627), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n776), .A2(new_n701), .A3(new_n750), .A4(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G122), .ZN(G24));
  NAND2_X1  g593(.A1(new_n637), .A2(G472), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n780), .A2(new_n769), .B1(new_n432), .B2(new_n774), .ZN(new_n781));
  NAND4_X1  g595(.A1(new_n781), .A2(new_n710), .A3(new_n744), .A4(new_n772), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n762), .ZN(new_n783));
  XNOR2_X1  g597(.A(KEYINPUT108), .B(G125), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n783), .B(new_n784), .ZN(G27));
  AOI21_X1  g599(.A(KEYINPUT32), .B1(new_n451), .B2(new_n432), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n452), .B(new_n447), .C1(new_n786), .C2(KEYINPUT110), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT110), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n434), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n515), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g604(.A1(new_n190), .A2(new_n307), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n386), .A2(new_n388), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n293), .A2(KEYINPUT109), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT109), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n292), .A2(new_n794), .A3(new_n195), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n283), .A2(G469), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n295), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n792), .B(new_n744), .C1(new_n797), .C2(new_n304), .ZN(new_n798));
  OAI21_X1  g612(.A(KEYINPUT42), .B1(new_n790), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n792), .B1(new_n797), .B2(new_n304), .ZN(new_n800));
  INV_X1    g614(.A(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(new_n704), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n669), .A2(new_n670), .A3(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(KEYINPUT42), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n801), .A2(new_n748), .A3(new_n804), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n799), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G131), .ZN(G33));
  NAND2_X1  g621(.A1(new_n453), .A2(new_n515), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n800), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n705), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(G134), .ZN(G36));
  OR2_X1    g625(.A1(new_n716), .A2(KEYINPUT45), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n283), .A2(KEYINPUT45), .A3(new_n793), .A4(new_n795), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n812), .A2(G469), .A3(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n814), .A2(KEYINPUT46), .A3(new_n295), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT46), .B1(new_n814), .B2(new_n295), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n815), .A2(new_n816), .A3(new_n304), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n190), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n386), .A2(new_n306), .A3(new_n388), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n664), .A2(new_n670), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT43), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT111), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT43), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n820), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT111), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n686), .B1(new_n638), .B2(new_n642), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n823), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT44), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n819), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n823), .A2(new_n826), .A3(KEYINPUT44), .A4(new_n827), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n818), .A2(new_n830), .A3(new_n722), .A4(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(G137), .ZN(G39));
  INV_X1    g647(.A(KEYINPUT47), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n817), .B2(new_n190), .ZN(new_n835));
  OR2_X1    g649(.A1(new_n816), .A2(new_n304), .ZN(new_n836));
  OAI211_X1 g650(.A(KEYINPUT47), .B(new_n191), .C1(new_n836), .C2(new_n815), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NOR4_X1   g652(.A1(new_n453), .A2(new_n515), .A3(new_n803), .A4(new_n819), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT112), .Z(new_n840));
  NOR2_X1   g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(new_n459), .ZN(G42));
  NOR2_X1   g656(.A1(new_n825), .A2(new_n626), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n843), .A2(new_n701), .A3(new_n750), .A4(new_n776), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT116), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n821), .A2(new_n776), .A3(new_n702), .ZN(new_n846));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n847), .A3(new_n701), .A4(new_n750), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n625), .ZN(new_n850));
  INV_X1    g664(.A(new_n819), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n750), .A2(new_n851), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n735), .A2(new_n852), .A3(new_n514), .A4(new_n626), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n850), .B1(new_n853), .B2(new_n751), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT117), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n849), .A2(new_n854), .A3(KEYINPUT117), .ZN(new_n858));
  INV_X1    g672(.A(new_n852), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n843), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n790), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT48), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n857), .A2(new_n858), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT118), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n857), .A2(KEYINPUT118), .A3(new_n858), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n749), .A2(new_n304), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n190), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n835), .A2(new_n837), .A3(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n846), .A2(new_n851), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n736), .A2(new_n515), .A3(new_n702), .A4(new_n859), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n664), .A2(new_n631), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n781), .A2(new_n710), .A3(new_n772), .ZN(new_n876));
  OAI22_X1  g690(.A1(new_n874), .A2(new_n875), .B1(new_n860), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n739), .A2(new_n306), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n846), .A2(new_n750), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT50), .ZN(new_n880));
  OR2_X1    g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n880), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n877), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n873), .A2(KEYINPUT51), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT51), .B1(new_n873), .B2(new_n883), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n778), .A2(new_n753), .A3(new_n756), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n887), .A2(new_n806), .A3(new_n767), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT114), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n631), .A2(new_n617), .A3(new_n802), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n686), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n453), .A2(new_n851), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n889), .B1(new_n892), .B2(new_n305), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n819), .A2(new_n686), .A3(new_n890), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n721), .A2(KEYINPUT114), .A3(new_n894), .A4(new_n453), .ZN(new_n895));
  AOI22_X1  g709(.A1(new_n893), .A2(new_n895), .B1(new_n809), .B2(new_n705), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n664), .A2(new_n631), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n897), .A2(new_n389), .A3(new_n627), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT113), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n389), .A2(new_n676), .A3(new_n627), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n897), .A2(new_n389), .A3(KEYINPUT113), .A4(new_n627), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n900), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n644), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n391), .B1(new_n688), .B2(new_n634), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n771), .A2(new_n775), .ZN(new_n906));
  INV_X1    g720(.A(new_n772), .ZN(new_n907));
  NOR4_X1   g721(.A1(new_n906), .A2(new_n907), .A3(new_n686), .A4(new_n803), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n801), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n896), .A2(new_n904), .A3(new_n905), .A4(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n888), .A2(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(new_n762), .ZN(new_n912));
  INV_X1    g726(.A(new_n706), .ZN(new_n913));
  INV_X1    g727(.A(new_n711), .ZN(new_n914));
  AOI22_X1  g728(.A1(new_n908), .A2(new_n912), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n710), .A2(new_n190), .A3(new_n704), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n797), .B2(new_n304), .ZN(new_n917));
  INV_X1    g731(.A(new_n734), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n646), .A2(new_n647), .A3(new_n740), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  NOR2_X1   g734(.A1(new_n920), .A2(new_n746), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n915), .A2(new_n921), .A3(KEYINPUT52), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT52), .ZN(new_n923));
  OAI22_X1  g737(.A1(new_n782), .A2(new_n762), .B1(new_n711), .B2(new_n706), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n734), .B(new_n916), .C1(new_n304), .C2(new_n797), .ZN(new_n925));
  OAI22_X1  g739(.A1(new_n925), .A2(new_n919), .B1(new_n745), .B2(new_n711), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n923), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT53), .B1(new_n911), .B2(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n764), .A2(new_n766), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n778), .A2(new_n753), .A3(new_n756), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n799), .A2(new_n805), .ZN(new_n932));
  NOR3_X1   g746(.A1(new_n930), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n893), .A2(new_n895), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n934), .A2(new_n909), .A3(new_n810), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n904), .A2(new_n905), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  AND4_X1   g751(.A1(KEYINPUT53), .A2(new_n928), .A3(new_n933), .A4(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT54), .B1(new_n929), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n928), .A2(new_n933), .A3(new_n937), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT53), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT54), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n748), .B(new_n750), .C1(new_n672), .C2(new_n677), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n767), .A2(new_n778), .A3(new_n944), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT115), .B1(new_n945), .B2(new_n932), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n935), .A2(new_n936), .A3(new_n941), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT115), .ZN(new_n948));
  NAND4_X1  g762(.A1(new_n887), .A2(new_n806), .A3(new_n948), .A4(new_n767), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n946), .A2(new_n947), .A3(new_n928), .A4(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n942), .A2(new_n943), .A3(new_n950), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n868), .A2(new_n886), .A3(new_n939), .A4(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(G952), .A2(G953), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT119), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT49), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n869), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT49), .B1(new_n749), .B2(new_n304), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n515), .A2(new_n820), .A3(new_n791), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n739), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n736), .A2(new_n957), .A3(new_n958), .A4(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n955), .A2(new_n961), .ZN(G75));
  INV_X1    g776(.A(KEYINPUT121), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n193), .A2(G952), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n189), .B(new_n387), .C1(new_n942), .C2(new_n950), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n346), .B(new_n360), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT55), .ZN(new_n968));
  XNOR2_X1  g782(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n965), .B1(new_n966), .B2(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(new_n968), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n942), .A2(new_n950), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(G902), .A3(new_n385), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT56), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n963), .B1(new_n972), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n968), .B1(new_n966), .B2(KEYINPUT56), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n964), .B1(new_n975), .B2(new_n970), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n979), .A2(new_n980), .A3(KEYINPUT121), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n978), .A2(new_n981), .ZN(G51));
  AOI21_X1  g796(.A(new_n189), .B1(new_n942), .B2(new_n950), .ZN(new_n983));
  INV_X1    g797(.A(new_n814), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n983), .A2(KEYINPUT122), .A3(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(KEYINPUT122), .B1(new_n983), .B2(new_n984), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n295), .B(KEYINPUT57), .Z(new_n988));
  AND3_X1   g802(.A1(new_n942), .A2(new_n943), .A3(new_n950), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n943), .B1(new_n942), .B2(new_n950), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n718), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n964), .B1(new_n987), .B2(new_n992), .ZN(G54));
  NOR2_X1   g807(.A1(new_n564), .A2(new_n544), .ZN(new_n994));
  INV_X1    g808(.A(new_n983), .ZN(new_n995));
  NAND2_X1  g809(.A1(KEYINPUT58), .A2(G475), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n965), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n995), .A2(new_n994), .A3(new_n996), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n998), .A2(new_n999), .ZN(G60));
  NAND2_X1  g814(.A1(G478), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT59), .Z(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(new_n939), .B2(new_n951), .ZN(new_n1003));
  OAI21_X1  g817(.A(KEYINPUT123), .B1(new_n1003), .B2(new_n662), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1002), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n911), .A2(KEYINPUT53), .A3(new_n928), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n943), .B1(new_n942), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1005), .B1(new_n989), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT123), .ZN(new_n1009));
  INV_X1    g823(.A(new_n662), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n974), .A2(KEYINPUT54), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n951), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n1010), .A2(new_n1002), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n964), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AND3_X1   g829(.A1(new_n1004), .A2(new_n1011), .A3(new_n1015), .ZN(G63));
  NAND2_X1  g830(.A1(G217), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT60), .Z(new_n1018));
  NAND2_X1  g832(.A1(new_n974), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n497), .A2(new_n500), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n974), .A2(new_n684), .A3(new_n1018), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1021), .A2(new_n965), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT61), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g839(.A1(new_n1021), .A2(KEYINPUT61), .A3(new_n965), .A4(new_n1022), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(G66));
  INV_X1    g841(.A(new_n620), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n193), .B1(new_n1028), .B2(G224), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n945), .A2(new_n936), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1030), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1029), .B1(new_n1031), .B2(new_n193), .ZN(new_n1032));
  INV_X1    g846(.A(new_n346), .ZN(new_n1033));
  OAI21_X1  g847(.A(new_n1033), .B1(G898), .B2(new_n193), .ZN(new_n1034));
  XOR2_X1   g848(.A(new_n1032), .B(new_n1034), .Z(G69));
  AOI21_X1  g849(.A(new_n193), .B1(G227), .B2(G900), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n402), .A2(new_n409), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT124), .Z(new_n1038));
  XNOR2_X1  g852(.A(new_n1038), .B(new_n561), .ZN(new_n1039));
  XOR2_X1   g853(.A(new_n1039), .B(KEYINPUT125), .Z(new_n1040));
  INV_X1    g854(.A(KEYINPUT62), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n924), .A2(new_n746), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1042), .ZN(new_n1043));
  OR3_X1    g857(.A1(new_n742), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g858(.A(new_n1041), .B1(new_n742), .B2(new_n1043), .ZN(new_n1045));
  NAND2_X1  g859(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  OR2_X1    g860(.A1(new_n838), .A2(new_n840), .ZN(new_n1047));
  OAI21_X1  g861(.A(new_n851), .B1(new_n897), .B2(new_n676), .ZN(new_n1048));
  OR3_X1    g862(.A1(new_n723), .A2(new_n808), .A3(new_n1048), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n832), .A2(KEYINPUT126), .A3(new_n1049), .ZN(new_n1050));
  INV_X1    g864(.A(new_n1050), .ZN(new_n1051));
  AOI21_X1  g865(.A(KEYINPUT126), .B1(new_n832), .B2(new_n1049), .ZN(new_n1052));
  OAI211_X1 g866(.A(new_n1046), .B(new_n1047), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1040), .B1(new_n1053), .B2(new_n193), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n1039), .B1(G900), .B2(G953), .ZN(new_n1055));
  INV_X1    g869(.A(new_n1055), .ZN(new_n1056));
  NOR2_X1   g870(.A1(new_n790), .A2(new_n919), .ZN(new_n1057));
  NAND3_X1  g871(.A1(new_n818), .A2(new_n722), .A3(new_n1057), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n932), .B1(new_n705), .B2(new_n809), .ZN(new_n1059));
  NAND4_X1  g873(.A1(new_n832), .A2(new_n1058), .A3(new_n1059), .A4(new_n1042), .ZN(new_n1060));
  NOR2_X1   g874(.A1(new_n841), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n1056), .B1(new_n1061), .B2(new_n193), .ZN(new_n1062));
  OAI21_X1  g876(.A(new_n1036), .B1(new_n1054), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g877(.A(new_n1036), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n1061), .A2(new_n193), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n1065), .A2(new_n1055), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n832), .A2(new_n1049), .ZN(new_n1067));
  INV_X1    g881(.A(KEYINPUT126), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g883(.A(new_n841), .B1(new_n1069), .B2(new_n1050), .ZN(new_n1070));
  AOI21_X1  g884(.A(G953), .B1(new_n1070), .B2(new_n1046), .ZN(new_n1071));
  OAI211_X1 g885(.A(new_n1064), .B(new_n1066), .C1(new_n1071), .C2(new_n1040), .ZN(new_n1072));
  NAND2_X1  g886(.A1(new_n1063), .A2(new_n1072), .ZN(G72));
  XNOR2_X1  g887(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1074));
  NOR2_X1   g888(.A1(new_n770), .A2(new_n189), .ZN(new_n1075));
  XOR2_X1   g889(.A(new_n1074), .B(new_n1075), .Z(new_n1076));
  INV_X1    g890(.A(new_n1076), .ZN(new_n1077));
  NOR2_X1   g891(.A1(new_n410), .A2(new_n418), .ZN(new_n1078));
  OAI221_X1 g892(.A(new_n1077), .B1(new_n1078), .B2(new_n438), .C1(new_n929), .C2(new_n938), .ZN(new_n1079));
  AOI21_X1  g893(.A(new_n1076), .B1(new_n1061), .B2(new_n1030), .ZN(new_n1080));
  NAND3_X1  g894(.A1(new_n421), .A2(new_n412), .A3(new_n430), .ZN(new_n1081));
  OAI211_X1 g895(.A(new_n965), .B(new_n1079), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g896(.A(new_n1077), .B1(new_n1053), .B2(new_n1031), .ZN(new_n1083));
  AOI21_X1  g897(.A(new_n1082), .B1(new_n730), .B2(new_n1083), .ZN(G57));
endmodule


