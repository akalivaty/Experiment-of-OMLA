//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1190, new_n1191, new_n1192, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n207));
  INV_X1    g0007(.A(G68), .ZN(new_n208));
  INV_X1    g0008(.A(G238), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n206), .B(new_n207), .C1(new_n208), .C2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT64), .ZN(new_n212));
  AOI211_X1 g0012(.A(new_n210), .B(new_n212), .C1(G77), .C2(G244), .ZN(new_n213));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n213), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT1), .Z(new_n218));
  OAI21_X1  g0018(.A(G50), .B1(G58), .B2(G68), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  NOR3_X1   g0020(.A1(new_n219), .A2(new_n215), .A3(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G13), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT0), .Z(new_n226));
  NOR3_X1   g0026(.A1(new_n218), .A2(new_n221), .A3(new_n226), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(G250), .B(G257), .Z(new_n232));
  XNOR2_X1  g0032(.A(G264), .B(G270), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n231), .B(new_n234), .ZN(G358));
  XNOR2_X1  g0035(.A(G68), .B(G77), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G50), .B(G58), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G87), .B(G116), .ZN(new_n239));
  INV_X1    g0039(.A(G107), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G97), .ZN(new_n241));
  INV_X1    g0041(.A(G97), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G107), .ZN(new_n243));
  NAND3_X1  g0043(.A1(new_n239), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G97), .B(G107), .ZN(new_n245));
  OAI21_X1  g0045(.A(new_n244), .B1(new_n239), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n238), .B(new_n246), .ZN(G351));
  XOR2_X1   g0047(.A(KEYINPUT8), .B(G58), .Z(new_n248));
  INV_X1    g0048(.A(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G20), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n248), .A2(new_n250), .B1(G20), .B2(new_n203), .ZN(new_n251));
  INV_X1    g0051(.A(G150), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n251), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n220), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NOR3_X1   g0058(.A1(new_n222), .A2(new_n215), .A3(G1), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n202), .ZN(new_n261));
  INV_X1    g0061(.A(new_n257), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G1), .B2(new_n215), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n261), .B1(new_n264), .B2(new_n202), .ZN(new_n265));
  AND2_X1   g0065(.A1(new_n265), .A2(KEYINPUT67), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(KEYINPUT67), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n258), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  OR2_X1    g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT66), .B(G1698), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n273), .B1(G222), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G223), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  OAI21_X1  g0077(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G41), .ZN(new_n279));
  OAI211_X1 g0079(.A(G1), .B(G13), .C1(new_n249), .C2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  OR2_X1    g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  OAI211_X1 g0084(.A(new_n278), .B(new_n281), .C1(G77), .C2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n279), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G226), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n214), .B1(G41), .B2(G45), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n280), .B1(KEYINPUT65), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT65), .ZN(new_n292));
  OAI21_X1  g0092(.A(G274), .B1(new_n287), .B2(new_n292), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n285), .A2(new_n289), .A3(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(G200), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n268), .A2(new_n269), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n270), .A2(new_n296), .A3(new_n297), .A4(new_n299), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT10), .ZN(new_n301));
  OR2_X1    g0101(.A1(new_n295), .A2(G179), .ZN(new_n302));
  INV_X1    g0102(.A(G169), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n295), .A2(new_n303), .ZN(new_n304));
  AND3_X1   g0104(.A1(new_n302), .A2(new_n268), .A3(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(G232), .ZN(new_n310));
  OAI221_X1 g0110(.A(new_n284), .B1(new_n209), .B2(new_n277), .C1(new_n309), .C2(new_n310), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n311), .B(new_n281), .C1(G107), .C2(new_n284), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n288), .A2(G244), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(new_n294), .A3(new_n313), .ZN(new_n314));
  XOR2_X1   g0114(.A(new_n314), .B(KEYINPUT68), .Z(new_n315));
  NOR2_X1   g0115(.A1(new_n315), .A2(new_n298), .ZN(new_n316));
  XOR2_X1   g0116(.A(KEYINPUT15), .B(G87), .Z(new_n317));
  AOI22_X1  g0117(.A1(new_n253), .A2(new_n248), .B1(new_n317), .B2(new_n250), .ZN(new_n318));
  INV_X1    g0118(.A(G77), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n318), .B1(new_n215), .B2(new_n319), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n320), .A2(new_n257), .B1(new_n319), .B2(new_n259), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n264), .A2(G77), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n314), .B(KEYINPUT68), .ZN(new_n325));
  INV_X1    g0125(.A(G200), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n316), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n315), .A2(new_n303), .ZN(new_n329));
  INV_X1    g0129(.A(G179), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n329), .A2(new_n323), .A3(new_n331), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n328), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g0133(.A(new_n301), .B(new_n306), .C1(new_n333), .C2(KEYINPUT69), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n328), .A2(KEYINPUT69), .A3(new_n332), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT14), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n274), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(new_n273), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n249), .A2(new_n242), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n281), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n288), .A2(G238), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n294), .A3(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n342), .B(KEYINPUT13), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n336), .B1(new_n343), .B2(G169), .ZN(new_n344));
  INV_X1    g0144(.A(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(new_n343), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G179), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n343), .A2(new_n336), .A3(G169), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n250), .A2(G77), .B1(new_n253), .B2(G50), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n215), .B2(G68), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n257), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n352), .B(KEYINPUT11), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n264), .A2(G68), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT70), .B1(new_n259), .B2(new_n208), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT12), .ZN(new_n356));
  AND3_X1   g0156(.A1(new_n353), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n349), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n358), .B1(new_n346), .B2(G190), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n326), .B2(new_n346), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n335), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n282), .A2(new_n215), .A3(new_n283), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT7), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n215), .A4(new_n283), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n208), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G58), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n368), .A2(new_n208), .ZN(new_n369));
  OAI21_X1  g0169(.A(G20), .B1(new_n369), .B2(new_n201), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n253), .A2(G159), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT16), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(KEYINPUT7), .B1(new_n273), .B2(new_n215), .ZN(new_n374));
  NOR4_X1   g0174(.A1(new_n271), .A2(new_n272), .A3(new_n364), .A4(G20), .ZN(new_n375));
  OAI21_X1  g0175(.A(G68), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT16), .ZN(new_n377));
  INV_X1    g0177(.A(new_n372), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n380), .A3(new_n377), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n373), .A2(new_n379), .A3(new_n381), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n376), .A2(new_n380), .A3(new_n377), .A4(new_n378), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n382), .A2(new_n257), .A3(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n260), .A2(new_n248), .ZN(new_n385));
  AOI21_X1  g0185(.A(new_n385), .B1(new_n264), .B2(new_n248), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n291), .A2(new_n293), .ZN(new_n388));
  NAND2_X1  g0188(.A1(G33), .A2(G87), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G226), .A2(G1698), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n274), .B2(G223), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n389), .B1(new_n392), .B2(new_n273), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n388), .B1(new_n393), .B2(new_n281), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n288), .A2(G232), .ZN(new_n395));
  AOI21_X1  g0195(.A(G169), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(G223), .B1(new_n307), .B2(new_n308), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n273), .B1(new_n397), .B2(new_n390), .ZN(new_n398));
  INV_X1    g0198(.A(new_n389), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n281), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND4_X1  g0200(.A1(new_n400), .A2(new_n330), .A3(new_n294), .A4(new_n395), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(KEYINPUT72), .B1(new_n396), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n400), .A2(new_n294), .A3(new_n395), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n303), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT72), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n406), .A3(new_n401), .ZN(new_n407));
  NAND4_X1  g0207(.A1(new_n387), .A2(KEYINPUT18), .A3(new_n403), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT73), .ZN(new_n409));
  AND3_X1   g0209(.A1(new_n405), .A2(new_n406), .A3(new_n401), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n406), .B1(new_n405), .B2(new_n401), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT73), .ZN(new_n413));
  NAND4_X1  g0213(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT18), .A4(new_n387), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT18), .ZN(new_n415));
  INV_X1    g0215(.A(new_n387), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n403), .A2(new_n407), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n409), .A2(new_n414), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n394), .A2(G190), .A3(new_n395), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n404), .A2(G200), .ZN(new_n421));
  NAND4_X1  g0221(.A1(new_n384), .A2(new_n420), .A3(new_n421), .A4(new_n386), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n422), .B(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NOR3_X1   g0224(.A1(new_n334), .A2(new_n362), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n215), .A2(G33), .A3(G116), .ZN(new_n426));
  XOR2_X1   g0226(.A(new_n426), .B(KEYINPUT85), .Z(new_n427));
  NOR2_X1   g0227(.A1(new_n273), .A2(G20), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT22), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n428), .A2(KEYINPUT84), .A3(new_n429), .A4(G87), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n284), .A2(KEYINPUT84), .A3(new_n215), .A4(G87), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT22), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n427), .B1(new_n430), .B2(new_n432), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n215), .A2(G107), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT23), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT86), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT24), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n433), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n436), .A2(KEYINPUT24), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(new_n439), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n433), .A2(new_n435), .A3(new_n437), .A4(new_n441), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n257), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT75), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n249), .A2(G1), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n259), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n444), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n447), .A2(new_n257), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(G107), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n259), .A2(new_n240), .ZN(new_n452));
  XOR2_X1   g0252(.A(new_n452), .B(KEYINPUT25), .Z(new_n453));
  NAND3_X1  g0253(.A1(new_n443), .A2(new_n451), .A3(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n279), .A2(KEYINPUT5), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n279), .A2(KEYINPUT5), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n286), .A2(G1), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n455), .A2(G274), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(G257), .B(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G294), .ZN(new_n460));
  OAI21_X1  g0260(.A(G250), .B1(new_n271), .B2(new_n272), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n459), .B(new_n460), .C1(new_n461), .C2(new_n309), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n281), .ZN(new_n463));
  INV_X1    g0263(.A(new_n456), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n214), .B(G45), .C1(new_n279), .C2(KEYINPUT5), .ZN(new_n465));
  OAI211_X1 g0265(.A(G264), .B(new_n280), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  AND3_X1   g0266(.A1(new_n463), .A2(KEYINPUT88), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(KEYINPUT88), .B1(new_n463), .B2(new_n466), .ZN(new_n468));
  OAI211_X1 g0268(.A(G179), .B(new_n458), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G250), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n470), .B1(new_n282), .B2(new_n283), .ZN(new_n471));
  AOI22_X1  g0271(.A1(new_n471), .A2(new_n274), .B1(G33), .B2(G294), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n280), .B1(new_n472), .B2(new_n459), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n458), .B1(new_n473), .B2(KEYINPUT87), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT87), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n466), .B1(new_n463), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g0276(.A(G169), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT89), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n469), .A2(new_n477), .A3(KEYINPUT89), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n454), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n466), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n483), .B1(new_n473), .B2(KEYINPUT87), .ZN(new_n484));
  INV_X1    g0284(.A(new_n458), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n485), .B1(new_n463), .B2(new_n475), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n298), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT88), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n488), .B1(new_n473), .B2(new_n483), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n463), .A2(KEYINPUT88), .A3(new_n466), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n485), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n487), .B1(new_n491), .B2(G200), .ZN(new_n492));
  NAND4_X1  g0292(.A1(new_n492), .A2(new_n451), .A3(new_n443), .A4(new_n453), .ZN(new_n493));
  INV_X1    g0293(.A(new_n457), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n280), .A2(new_n494), .A3(G250), .ZN(new_n495));
  INV_X1    g0295(.A(G274), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(new_n494), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT76), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT76), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n495), .B(new_n499), .C1(new_n496), .C2(new_n494), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n274), .A2(G238), .B1(G244), .B2(G1698), .ZN(new_n502));
  INV_X1    g0302(.A(G116), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n502), .A2(new_n273), .B1(new_n249), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n281), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n428), .A2(G68), .ZN(new_n507));
  XOR2_X1   g0307(.A(KEYINPUT77), .B(KEYINPUT19), .Z(new_n508));
  NOR3_X1   g0308(.A1(new_n249), .A2(new_n242), .A3(G20), .ZN(new_n509));
  XOR2_X1   g0309(.A(KEYINPUT78), .B(G87), .Z(new_n510));
  NOR3_X1   g0310(.A1(new_n510), .A2(G97), .A3(G107), .ZN(new_n511));
  AOI21_X1  g0311(.A(G20), .B1(new_n508), .B2(new_n339), .ZN(new_n512));
  OAI221_X1 g0312(.A(new_n507), .B1(new_n508), .B2(new_n509), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n317), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n513), .A2(new_n257), .B1(new_n259), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n450), .A2(new_n317), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n330), .A2(new_n506), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n501), .A2(new_n505), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(new_n303), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n482), .A2(new_n493), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n260), .A2(G97), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n450), .A2(G97), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n240), .B1(new_n365), .B2(new_n366), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT6), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n245), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n241), .A2(new_n526), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n215), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n254), .A2(new_n319), .ZN(new_n531));
  NOR3_X1   g0331(.A1(new_n525), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n532), .A2(KEYINPUT74), .A3(new_n262), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT74), .ZN(new_n534));
  OAI21_X1  g0334(.A(G107), .B1(new_n374), .B2(new_n375), .ZN(new_n535));
  INV_X1    g0335(.A(new_n531), .ZN(new_n536));
  INV_X1    g0336(.A(new_n527), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(new_n528), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n535), .B(new_n536), .C1(new_n538), .C2(new_n215), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n534), .B1(new_n539), .B2(new_n257), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n523), .B(new_n524), .C1(new_n533), .C2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(G257), .B(new_n280), .C1(new_n464), .C2(new_n465), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT4), .ZN(new_n544));
  OAI21_X1  g0344(.A(G244), .B1(new_n307), .B2(new_n308), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n544), .B1(new_n545), .B2(new_n273), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n284), .A2(new_n274), .A3(KEYINPUT4), .A4(G244), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n471), .A2(G1698), .ZN(new_n548));
  NAND2_X1  g0348(.A1(G33), .A2(G283), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n546), .A2(new_n547), .A3(new_n548), .A4(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n543), .B1(new_n550), .B2(new_n281), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n551), .A2(new_n330), .A3(new_n458), .ZN(new_n552));
  AOI21_X1  g0352(.A(G169), .B1(new_n551), .B2(new_n458), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n541), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n450), .A2(G87), .ZN(new_n556));
  AND2_X1   g0356(.A1(new_n515), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n506), .A2(G190), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n518), .A2(G200), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n557), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(KEYINPUT74), .B1(new_n532), .B2(new_n262), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n539), .A2(new_n534), .A3(new_n257), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n522), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n551), .A2(new_n298), .A3(new_n458), .ZN(new_n564));
  AOI211_X1 g0364(.A(new_n543), .B(new_n485), .C1(new_n550), .C2(new_n281), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(G200), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n563), .A2(new_n566), .A3(new_n524), .ZN(new_n567));
  AND3_X1   g0367(.A1(new_n555), .A2(new_n560), .A3(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT21), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT80), .ZN(new_n570));
  OAI21_X1  g0370(.A(G257), .B1(new_n271), .B2(new_n272), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n570), .B1(new_n571), .B2(new_n309), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n284), .A2(new_n274), .A3(KEYINPUT80), .A4(G257), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n273), .A2(G303), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n284), .A2(G264), .A3(G1698), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n572), .A2(new_n573), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT81), .ZN(new_n577));
  AND3_X1   g0377(.A1(new_n576), .A2(new_n577), .A3(new_n281), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n577), .B1(new_n576), .B2(new_n281), .ZN(new_n579));
  OAI211_X1 g0379(.A(G270), .B(new_n280), .C1(new_n464), .C2(new_n465), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT79), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n580), .A2(new_n581), .A3(new_n458), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n581), .B1(new_n580), .B2(new_n458), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n578), .A2(new_n579), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n259), .A2(new_n503), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n549), .B(new_n215), .C1(G33), .C2(new_n242), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n587), .B(new_n257), .C1(new_n215), .C2(G116), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT20), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  OAI221_X1 g0391(.A(new_n586), .B1(new_n449), .B2(new_n503), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G169), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n569), .B1(new_n585), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT83), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT83), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n596), .B(new_n569), .C1(new_n585), .C2(new_n593), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n585), .A2(G179), .A3(new_n592), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n576), .A2(new_n281), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(KEYINPUT81), .ZN(new_n601));
  OR2_X1    g0401(.A1(new_n582), .A2(new_n583), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n576), .A2(new_n577), .A3(new_n281), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n601), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n604), .A2(KEYINPUT21), .A3(G169), .A4(new_n592), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n599), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(KEYINPUT82), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT82), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n599), .A2(new_n605), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(G200), .ZN(new_n610));
  INV_X1    g0410(.A(new_n592), .ZN(new_n611));
  OAI211_X1 g0411(.A(new_n610), .B(new_n611), .C1(new_n298), .C2(new_n604), .ZN(new_n612));
  AND4_X1   g0412(.A1(new_n598), .A2(new_n607), .A3(new_n609), .A4(new_n612), .ZN(new_n613));
  AND4_X1   g0413(.A1(new_n425), .A2(new_n521), .A3(new_n568), .A4(new_n613), .ZN(G372));
  NAND2_X1  g0414(.A1(new_n418), .A2(new_n408), .ZN(new_n615));
  INV_X1    g0415(.A(new_n348), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n344), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n357), .B1(new_n617), .B2(new_n347), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n329), .A2(new_n323), .A3(new_n331), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n619), .B2(new_n361), .ZN(new_n620));
  INV_X1    g0420(.A(new_n423), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n615), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n305), .B1(new_n622), .B2(new_n301), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT91), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n493), .A2(new_n555), .A3(new_n567), .A4(new_n560), .ZN(new_n625));
  AND2_X1   g0425(.A1(new_n519), .A2(KEYINPUT90), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n519), .A2(KEYINPUT90), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n517), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n624), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n568), .A2(KEYINPUT91), .A3(new_n493), .A4(new_n628), .ZN(new_n631));
  INV_X1    g0431(.A(new_n606), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n454), .A2(new_n478), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n598), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n630), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n520), .A2(new_n560), .A3(new_n541), .A4(new_n554), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(KEYINPUT26), .ZN(new_n637));
  INV_X1    g0437(.A(new_n555), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n638), .A2(new_n628), .A3(new_n639), .A4(new_n560), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n637), .A2(new_n640), .A3(new_n628), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n635), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n425), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n623), .A2(new_n643), .ZN(G369));
  NAND2_X1  g0444(.A1(new_n598), .A2(new_n632), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n222), .A2(G20), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n646), .A2(new_n214), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(KEYINPUT27), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n648), .A2(G213), .A3(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(G343), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n592), .A2(new_n652), .ZN(new_n653));
  MUX2_X1   g0453(.A(new_n645), .B(new_n613), .S(new_n653), .Z(new_n654));
  XOR2_X1   g0454(.A(new_n654), .B(KEYINPUT92), .Z(new_n655));
  AND2_X1   g0455(.A1(new_n655), .A2(G330), .ZN(new_n656));
  INV_X1    g0456(.A(new_n652), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n482), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n454), .A2(new_n652), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n482), .A2(new_n493), .A3(new_n659), .ZN(new_n660));
  AND3_X1   g0460(.A1(new_n658), .A2(KEYINPUT93), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(KEYINPUT93), .B1(new_n658), .B2(new_n660), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n656), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g0465(.A(new_n665), .B(KEYINPUT94), .Z(new_n666));
  AND3_X1   g0466(.A1(new_n598), .A2(new_n607), .A3(new_n609), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n667), .A2(new_n652), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n633), .A2(new_n652), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n666), .A2(new_n673), .ZN(G399));
  NOR2_X1   g0474(.A1(new_n223), .A2(G41), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G1), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n511), .A2(new_n503), .ZN(new_n678));
  OAI22_X1  g0478(.A1(new_n677), .A2(new_n678), .B1(new_n219), .B2(new_n676), .ZN(new_n679));
  XNOR2_X1  g0479(.A(new_n679), .B(KEYINPUT28), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n613), .A2(new_n521), .A3(new_n568), .A4(new_n657), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n604), .A2(new_n330), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n489), .A2(new_n490), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(new_n506), .A4(new_n565), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT95), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(KEYINPUT30), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n684), .A2(new_n686), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n491), .A2(new_n565), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT96), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n691), .A2(new_n518), .A3(new_n604), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n330), .B1(new_n689), .B2(new_n690), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n687), .B(new_n688), .C1(new_n692), .C2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n652), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n681), .A2(new_n695), .A3(KEYINPUT31), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT31), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n694), .A2(new_n697), .A3(new_n652), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(G330), .ZN(new_n700));
  AOI211_X1 g0500(.A(KEYINPUT29), .B(new_n652), .C1(new_n635), .C2(new_n641), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n598), .A2(new_n482), .A3(new_n607), .A4(new_n609), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(new_n493), .A3(new_n568), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n638), .A2(new_n628), .A3(new_n560), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n629), .B1(new_n705), .B2(KEYINPUT26), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n636), .A2(KEYINPUT26), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n702), .B1(new_n708), .B2(new_n657), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n701), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n700), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n680), .B1(new_n712), .B2(G1), .ZN(G364));
  NOR2_X1   g0513(.A1(new_n219), .A2(G45), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n238), .A2(G45), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(KEYINPUT97), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n223), .A2(new_n284), .ZN(new_n717));
  OAI211_X1 g0517(.A(new_n716), .B(new_n717), .C1(KEYINPUT97), .C2(new_n715), .ZN(new_n718));
  INV_X1    g0518(.A(G355), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n224), .A2(new_n284), .ZN(new_n720));
  OAI221_X1 g0520(.A(new_n718), .B1(G116), .B2(new_n224), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(G13), .A2(G33), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G20), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n220), .B1(G20), .B2(new_n303), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n721), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n677), .B1(G45), .B2(new_n646), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n330), .A2(new_n326), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n215), .A2(G190), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(G317), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n733), .A2(KEYINPUT33), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n733), .A2(KEYINPUT33), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n732), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n215), .A2(new_n298), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n326), .A2(G179), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G303), .ZN(new_n740));
  INV_X1    g0540(.A(G322), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n330), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n737), .A2(new_n742), .ZN(new_n743));
  OAI221_X1 g0543(.A(new_n273), .B1(new_n739), .B2(new_n740), .C1(new_n741), .C2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G179), .A2(G200), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n215), .B1(new_n745), .B2(G190), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI211_X1 g0547(.A(new_n736), .B(new_n744), .C1(G294), .C2(new_n747), .ZN(new_n748));
  XNOR2_X1  g0548(.A(KEYINPUT98), .B(G326), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n730), .A2(new_n737), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n731), .A2(new_n742), .ZN(new_n752));
  INV_X1    g0552(.A(G311), .ZN(new_n753));
  OAI22_X1  g0553(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n731), .A2(new_n745), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n754), .B1(G329), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(G283), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n731), .A2(new_n738), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n748), .B(new_n757), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  XNOR2_X1  g0560(.A(new_n760), .B(KEYINPUT99), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n732), .A2(new_n208), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n756), .A2(G159), .ZN(new_n763));
  XNOR2_X1  g0563(.A(new_n763), .B(KEYINPUT32), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n746), .A2(new_n242), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n743), .A2(new_n368), .B1(new_n752), .B2(new_n319), .ZN(new_n767));
  INV_X1    g0567(.A(new_n739), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(new_n510), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n284), .B1(new_n751), .B2(new_n202), .ZN(new_n770));
  INV_X1    g0570(.A(new_n759), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n770), .B1(G107), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n766), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n761), .B1(new_n762), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n729), .B1(new_n774), .B2(new_n725), .ZN(new_n775));
  INV_X1    g0575(.A(new_n724), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n727), .B(new_n775), .C1(new_n654), .C2(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n655), .A2(G330), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n729), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n655), .A2(G330), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n777), .B1(new_n779), .B2(new_n780), .ZN(G396));
  AOI21_X1  g0581(.A(new_n652), .B1(new_n635), .B2(new_n641), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n619), .A2(new_n657), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n323), .A2(new_n652), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n784), .B1(new_n316), .B2(new_n327), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(new_n332), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n782), .A2(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n652), .B(new_n787), .C1(new_n635), .C2(new_n641), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(new_n700), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(new_n729), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n771), .A2(G87), .ZN(new_n794));
  INV_X1    g0594(.A(G294), .ZN(new_n795));
  OAI221_X1 g0595(.A(new_n794), .B1(new_n240), .B2(new_n739), .C1(new_n795), .C2(new_n743), .ZN(new_n796));
  INV_X1    g0596(.A(new_n752), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n796), .B1(G116), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n273), .B1(new_n732), .B2(new_n758), .ZN(new_n799));
  INV_X1    g0599(.A(new_n751), .ZN(new_n800));
  AOI211_X1 g0600(.A(new_n765), .B(new_n799), .C1(G303), .C2(new_n800), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n798), .B(new_n801), .C1(new_n753), .C2(new_n755), .ZN(new_n802));
  INV_X1    g0602(.A(new_n743), .ZN(new_n803));
  INV_X1    g0603(.A(new_n732), .ZN(new_n804));
  AOI22_X1  g0604(.A1(G143), .A2(new_n803), .B1(new_n804), .B2(G150), .ZN(new_n805));
  INV_X1    g0605(.A(G137), .ZN(new_n806));
  INV_X1    g0606(.A(G159), .ZN(new_n807));
  OAI221_X1 g0607(.A(new_n805), .B1(new_n806), .B2(new_n751), .C1(new_n807), .C2(new_n752), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT34), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n759), .A2(new_n208), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n284), .B1(new_n739), .B2(new_n202), .ZN(new_n813));
  AOI211_X1 g0613(.A(new_n812), .B(new_n813), .C1(G58), .C2(new_n747), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n810), .A2(new_n811), .A3(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n755), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n802), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n725), .A2(new_n722), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n818), .A2(new_n725), .B1(new_n319), .B2(new_n819), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n728), .B(new_n820), .C1(new_n788), .C2(new_n723), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n793), .A2(new_n821), .ZN(G384));
  AND2_X1   g0622(.A1(new_n373), .A2(new_n379), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n386), .B1(new_n823), .B2(new_n262), .ZN(new_n824));
  INV_X1    g0624(.A(new_n650), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n424), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT37), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n825), .B1(new_n403), .B2(new_n407), .ZN(new_n830));
  OAI211_X1 g0630(.A(new_n829), .B(new_n422), .C1(new_n830), .C2(new_n416), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n650), .B1(new_n410), .B2(new_n411), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n824), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n829), .B1(new_n834), .B2(new_n422), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n828), .A2(KEYINPUT38), .A3(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT39), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT38), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n833), .A2(new_n387), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(new_n422), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT101), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n833), .B2(new_n387), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n841), .B1(new_n829), .B2(new_n843), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n840), .A2(new_n842), .A3(KEYINPUT37), .A4(new_n422), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n387), .A2(new_n825), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n847), .B1(new_n615), .B2(new_n423), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n839), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n837), .A2(new_n838), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n826), .B1(new_n419), .B2(new_n423), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n832), .A2(new_n835), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n839), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n838), .B1(new_n837), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g0654(.A(KEYINPUT102), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n359), .A2(new_n652), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT38), .B1(new_n828), .B2(new_n836), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n851), .A2(new_n852), .A3(new_n839), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT39), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT102), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n837), .A2(new_n838), .A3(new_n849), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n855), .A2(new_n856), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n615), .A2(new_n825), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n783), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n782), .B2(new_n788), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n857), .A2(new_n858), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT100), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n359), .B2(new_n657), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n618), .A2(KEYINPUT100), .A3(new_n652), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n359), .A2(new_n361), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n358), .A2(new_n652), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n870), .A2(new_n871), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OR3_X1    g0674(.A1(new_n867), .A2(new_n868), .A3(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n863), .A2(new_n865), .A3(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT103), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n863), .A2(new_n875), .A3(KEYINPUT103), .A4(new_n865), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n425), .B1(new_n701), .B2(new_n709), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n623), .ZN(new_n882));
  XOR2_X1   g0682(.A(new_n882), .B(KEYINPUT104), .Z(new_n883));
  XNOR2_X1  g0683(.A(new_n880), .B(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n359), .A2(new_n361), .A3(new_n873), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT100), .B1(new_n618), .B2(new_n652), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n359), .A2(new_n869), .A3(new_n657), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND4_X1  g0688(.A1(new_n888), .A2(new_n696), .A3(new_n698), .A4(new_n788), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n837), .A2(new_n849), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT40), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n889), .B2(new_n868), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n699), .A2(new_n425), .ZN(new_n896));
  XOR2_X1   g0696(.A(new_n895), .B(new_n896), .Z(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(G330), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n884), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n884), .A2(new_n898), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n899), .B1(KEYINPUT105), .B2(new_n900), .ZN(new_n901));
  OAI221_X1 g0701(.A(new_n901), .B1(KEYINPUT105), .B2(new_n900), .C1(new_n214), .C2(new_n646), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT35), .ZN(new_n903));
  AOI211_X1 g0703(.A(new_n215), .B(new_n220), .C1(new_n538), .C2(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n904), .B(G116), .C1(new_n903), .C2(new_n538), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT36), .ZN(new_n906));
  OAI21_X1  g0706(.A(G77), .B1(new_n368), .B2(new_n208), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n907), .A2(new_n219), .B1(G50), .B2(new_n208), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(G1), .A3(new_n222), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n902), .A2(new_n906), .A3(new_n909), .ZN(G367));
  NAND2_X1  g0710(.A1(new_n638), .A2(new_n652), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n541), .A2(new_n652), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n555), .A2(new_n912), .A3(new_n567), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n666), .A2(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(new_n628), .B(new_n560), .C1(new_n557), .C2(new_n657), .ZN(new_n917));
  OR2_X1    g0717(.A1(new_n917), .A2(KEYINPUT106), .ZN(new_n918));
  OR3_X1    g0718(.A1(new_n628), .A2(new_n557), .A3(new_n657), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(KEYINPUT106), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  XOR2_X1   g0721(.A(KEYINPUT107), .B(KEYINPUT43), .Z(new_n922));
  NOR2_X1   g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n664), .A2(new_n668), .A3(new_n914), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT42), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n924), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n555), .B1(new_n913), .B2(new_n482), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n657), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n923), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n926), .A2(new_n923), .A3(new_n928), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n916), .B(new_n933), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n675), .B(KEYINPUT41), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n665), .B(KEYINPUT94), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n672), .A2(new_n915), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT45), .ZN(new_n939));
  OAI211_X1 g0739(.A(KEYINPUT108), .B(KEYINPUT44), .C1(new_n673), .C2(new_n914), .ZN(new_n940));
  NAND2_X1  g0740(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n941));
  OR2_X1    g0741(.A1(KEYINPUT108), .A2(KEYINPUT44), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n672), .A2(new_n915), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n939), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n937), .A2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n937), .A2(new_n944), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n663), .B(new_n668), .Z(new_n948));
  XNOR2_X1  g0748(.A(new_n778), .B(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n949), .A2(new_n711), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n946), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n936), .B1(new_n951), .B2(new_n712), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n214), .B1(new_n646), .B2(G45), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT109), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n934), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n717), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n726), .B1(new_n224), .B2(new_n514), .C1(new_n234), .C2(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n755), .A2(new_n806), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n743), .A2(new_n252), .B1(new_n759), .B2(new_n319), .ZN(new_n959));
  AOI211_X1 g0759(.A(new_n958), .B(new_n959), .C1(G143), .C2(new_n800), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n746), .A2(new_n208), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n284), .B1(new_n739), .B2(new_n368), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n961), .B(new_n962), .C1(G50), .C2(new_n797), .ZN(new_n963));
  OAI211_X1 g0763(.A(new_n960), .B(new_n963), .C1(new_n807), .C2(new_n732), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n752), .A2(new_n758), .B1(new_n746), .B2(new_n240), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT110), .Z(new_n966));
  NOR2_X1   g0766(.A1(new_n759), .A2(new_n242), .ZN(new_n967));
  OAI22_X1  g0767(.A1(new_n743), .A2(new_n740), .B1(new_n755), .B2(new_n733), .ZN(new_n968));
  AOI211_X1 g0768(.A(new_n967), .B(new_n968), .C1(G294), .C2(new_n804), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n768), .A2(KEYINPUT46), .A3(G116), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT46), .B1(new_n768), .B2(G116), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n971), .A2(new_n284), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n966), .A2(new_n969), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n751), .A2(new_n753), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n964), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XNOR2_X1  g0775(.A(new_n975), .B(KEYINPUT47), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n729), .B1(new_n976), .B2(new_n725), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n957), .B(new_n977), .C1(new_n921), .C2(new_n776), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n955), .A2(new_n978), .ZN(G387));
  OR3_X1    g0779(.A1(new_n950), .A2(KEYINPUT112), .A3(new_n676), .ZN(new_n980));
  OAI21_X1  g0780(.A(KEYINPUT112), .B1(new_n950), .B2(new_n676), .ZN(new_n981));
  INV_X1    g0781(.A(new_n949), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n980), .B(new_n981), .C1(new_n712), .C2(new_n982), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n954), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n273), .B1(new_n759), .B2(new_n503), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G311), .A2(new_n804), .B1(new_n803), .B2(G317), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n740), .B2(new_n752), .C1(new_n741), .C2(new_n751), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT48), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n758), .B2(new_n746), .C1(new_n795), .C2(new_n739), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT49), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n985), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n990), .B2(new_n989), .C1(new_n755), .C2(new_n750), .ZN(new_n992));
  INV_X1    g0792(.A(new_n248), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(new_n732), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n768), .A2(G77), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n995), .B1(new_n755), .B2(new_n252), .C1(new_n208), .C2(new_n752), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G159), .B2(new_n800), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n747), .A2(new_n317), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n273), .B(new_n967), .C1(G50), .C2(new_n803), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n992), .B1(new_n994), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n717), .B1(new_n231), .B2(new_n286), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n678), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1002), .B1(new_n1003), .B2(new_n720), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n1003), .B(new_n286), .C1(new_n208), .C2(new_n319), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n248), .A2(new_n202), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1006), .B(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1004), .B1(new_n1005), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(G107), .B2(new_n224), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1001), .A2(new_n725), .B1(new_n726), .B2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n1011), .B(new_n728), .C1(new_n664), .C2(new_n776), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n983), .A2(new_n984), .A3(new_n1012), .ZN(G393));
  OAI22_X1  g0813(.A1(new_n751), .A2(new_n733), .B1(new_n743), .B2(new_n753), .ZN(new_n1014));
  XOR2_X1   g0814(.A(new_n1014), .B(KEYINPUT114), .Z(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT52), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(G294), .A2(new_n797), .B1(new_n756), .B2(G322), .ZN(new_n1017));
  OAI221_X1 g0817(.A(new_n1017), .B1(new_n758), .B2(new_n739), .C1(new_n740), .C2(new_n732), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G107), .B2(new_n771), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n284), .B1(new_n747), .B2(G116), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1016), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G68), .A2(new_n768), .B1(new_n756), .B2(G143), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n1022), .B1(new_n202), .B2(new_n732), .C1(new_n993), .C2(new_n752), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(G77), .B2(new_n747), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n751), .A2(new_n252), .B1(new_n743), .B2(new_n807), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT51), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1024), .A2(new_n284), .A3(new_n794), .A4(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1021), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n725), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n246), .A2(new_n717), .B1(G97), .B2(new_n223), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n729), .B1(new_n1030), .B2(new_n726), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT113), .Z(new_n1032));
  OAI211_X1 g0832(.A(new_n1029), .B(new_n1032), .C1(new_n914), .C2(new_n776), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n950), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n947), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1035), .B1(new_n1036), .B2(new_n945), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n1037), .A2(new_n951), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1034), .B1(new_n1038), .B2(new_n675), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n946), .A2(new_n947), .A3(new_n954), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(G390));
  NAND4_X1  g0841(.A1(new_n696), .A2(G330), .A3(new_n698), .A4(new_n788), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1042), .A2(new_n874), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n888), .B1(new_n790), .B2(new_n866), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n856), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n855), .A2(new_n862), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n890), .A2(new_n1045), .ZN(new_n1047));
  AND2_X1   g0847(.A1(new_n708), .A2(new_n657), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n786), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n783), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1047), .B1(new_n1050), .B2(new_n888), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1043), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1045), .B1(new_n867), .B2(new_n874), .ZN(new_n1053));
  NOR3_X1   g0853(.A1(new_n850), .A2(new_n854), .A3(KEYINPUT102), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n860), .B1(new_n859), .B2(new_n861), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1053), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n866), .B1(new_n1048), .B2(new_n786), .ZN(new_n1057));
  OAI211_X1 g0857(.A(new_n1045), .B(new_n890), .C1(new_n1057), .C2(new_n874), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n699), .A2(G330), .A3(new_n788), .A4(new_n888), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1052), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n954), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n722), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n751), .A2(new_n758), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n743), .A2(new_n503), .B1(new_n755), .B2(new_n795), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1065), .B(new_n1066), .C1(G87), .C2(new_n768), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n747), .A2(G77), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n797), .A2(G97), .ZN(new_n1069));
  AOI211_X1 g0869(.A(new_n284), .B(new_n812), .C1(G107), .C2(new_n804), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n739), .A2(new_n252), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT53), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n1072), .A2(new_n1073), .B1(new_n807), .B2(new_n746), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1072), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n284), .B1(new_n1075), .B2(KEYINPUT53), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n1074), .B(new_n1076), .C1(G50), .C2(new_n771), .ZN(new_n1077));
  INV_X1    g0877(.A(G128), .ZN(new_n1078));
  INV_X1    g0878(.A(G125), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n751), .A2(new_n1078), .B1(new_n755), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT115), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(KEYINPUT54), .B(G143), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n732), .A2(new_n806), .B1(new_n752), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1080), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1077), .B(new_n1084), .C1(new_n1081), .C2(new_n1083), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n743), .A2(new_n816), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1071), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1087), .A2(new_n725), .B1(new_n993), .B2(new_n819), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1064), .A2(new_n728), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n699), .A2(G330), .A3(new_n425), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n881), .A3(new_n623), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n867), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1042), .A2(new_n874), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1092), .B1(new_n1093), .B2(new_n1043), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1042), .A2(new_n874), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1059), .A2(new_n1057), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1091), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n1062), .A2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1052), .A2(new_n1097), .A3(new_n1060), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n675), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1063), .B(new_n1089), .C1(new_n1098), .C2(new_n1100), .ZN(G378));
  INV_X1    g0901(.A(KEYINPUT57), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1091), .ZN(new_n1103));
  AND3_X1   g0903(.A1(new_n1099), .A2(KEYINPUT119), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(KEYINPUT119), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n892), .A2(new_n894), .A3(G330), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n301), .A2(new_n306), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT55), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n268), .A2(new_n825), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT56), .Z(new_n1111));
  XNOR2_X1  g0911(.A(new_n1109), .B(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1107), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1112), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1114), .A2(new_n892), .A3(new_n894), .A4(G330), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n880), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g0917(.A1(new_n878), .A2(new_n1113), .A3(new_n879), .A4(new_n1115), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1102), .B1(new_n1106), .B2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1117), .A2(KEYINPUT57), .A3(new_n1118), .ZN(new_n1121));
  OAI21_X1  g0921(.A(KEYINPUT120), .B1(new_n1106), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1121), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT119), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1099), .A2(KEYINPUT119), .A3(new_n1103), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT120), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1123), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1120), .A2(new_n1122), .A3(new_n1130), .A4(new_n675), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1112), .A2(new_n722), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n202), .B1(new_n271), .B2(G41), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n732), .A2(new_n816), .B1(new_n752), .B2(new_n806), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT116), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n751), .A2(new_n1079), .B1(new_n739), .B2(new_n1082), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G150), .B2(new_n747), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(new_n1078), .C2(new_n743), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT59), .ZN(new_n1139));
  AOI21_X1  g0939(.A(G41), .B1(new_n756), .B2(G124), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1140), .B(new_n249), .C1(new_n807), .C2(new_n759), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT117), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1133), .B1(new_n1139), .B2(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(G116), .A2(new_n800), .B1(new_n804), .B2(G97), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n1144), .B1(new_n368), .B2(new_n759), .C1(new_n758), .C2(new_n755), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(G107), .A2(new_n803), .B1(new_n797), .B2(new_n317), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n961), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1146), .A2(new_n279), .A3(new_n1147), .A4(new_n995), .ZN(new_n1148));
  NOR3_X1   g0948(.A1(new_n1145), .A2(new_n284), .A3(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n1149), .B(KEYINPUT58), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n725), .B1(new_n1143), .B2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT118), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n202), .B2(new_n819), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1132), .A2(new_n728), .A3(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1119), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1156), .B2(new_n954), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1131), .A2(new_n1157), .ZN(G375));
  INV_X1    g0958(.A(new_n1097), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1094), .A2(new_n1091), .A3(new_n1096), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1159), .A2(new_n935), .A3(new_n1160), .ZN(new_n1161));
  XOR2_X1   g0961(.A(new_n954), .B(KEYINPUT121), .Z(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n874), .A2(new_n722), .ZN(new_n1165));
  OAI22_X1  g0965(.A1(new_n752), .A2(new_n252), .B1(new_n746), .B2(new_n202), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT123), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n732), .A2(new_n1082), .B1(new_n755), .B2(new_n1078), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n284), .B1(new_n759), .B2(new_n368), .C1(new_n806), .C2(new_n743), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n739), .A2(new_n807), .ZN(new_n1171));
  NOR4_X1   g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n1167), .B2(new_n1166), .C1(new_n816), .C2(new_n751), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n998), .B1(new_n758), .B2(new_n743), .ZN(new_n1174));
  XOR2_X1   g0974(.A(new_n1174), .B(KEYINPUT122), .Z(new_n1175));
  OAI22_X1  g0975(.A1(new_n751), .A2(new_n795), .B1(new_n739), .B2(new_n242), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n273), .B1(new_n755), .B2(new_n740), .C1(new_n319), .C2(new_n759), .ZN(new_n1177));
  AOI211_X1 g0977(.A(new_n1176), .B(new_n1177), .C1(G116), .C2(new_n804), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1175), .B(new_n1178), .C1(new_n240), .C2(new_n752), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1173), .A2(new_n1179), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(new_n1180), .A2(new_n725), .B1(new_n208), .B2(new_n819), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1165), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1164), .B1(new_n728), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1161), .A2(new_n1183), .ZN(G381));
  NAND4_X1  g0984(.A1(new_n1039), .A2(new_n955), .A3(new_n978), .A4(new_n1040), .ZN(new_n1185));
  OR2_X1    g0985(.A1(G393), .A2(G396), .ZN(new_n1186));
  NOR4_X1   g0986(.A1(new_n1185), .A2(G384), .A3(G381), .A4(new_n1186), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(G375), .A2(G378), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(G407));
  NAND2_X1  g0989(.A1(new_n651), .A2(G213), .ZN(new_n1190));
  XOR2_X1   g0990(.A(new_n1190), .B(KEYINPUT124), .Z(new_n1191));
  OAI21_X1  g0991(.A(new_n1188), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1192), .A2(G213), .ZN(G409));
  INV_X1    g0993(.A(KEYINPUT126), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1163), .B1(new_n1106), .B2(new_n936), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n1156), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G378), .B1(new_n1196), .B2(new_n1154), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1122), .A2(new_n1130), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1119), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n675), .B1(new_n1199), .B2(KEYINPUT57), .ZN(new_n1200));
  OAI211_X1 g1000(.A(G378), .B(new_n1157), .C1(new_n1198), .C2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(KEYINPUT125), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT125), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1131), .A2(new_n1203), .A3(G378), .A4(new_n1157), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1197), .B1(new_n1202), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(KEYINPUT60), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1160), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1160), .A2(new_n1206), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1207), .A2(new_n675), .A3(new_n1159), .A4(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1183), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(new_n793), .A3(new_n821), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1209), .A2(G384), .A3(new_n1183), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1205), .A2(new_n1191), .A3(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1191), .A2(G2897), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1213), .B(new_n1215), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1216), .B1(new_n1205), .B2(new_n1191), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1214), .B1(new_n1217), .B2(KEYINPUT63), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(G390), .A2(G387), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G393), .A2(G396), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1186), .A2(new_n1220), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1219), .A2(new_n1185), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1221), .B1(new_n1219), .B2(new_n1185), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1202), .A2(new_n1204), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1197), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1191), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1213), .ZN(new_n1229));
  NAND4_X1  g1029(.A1(new_n1227), .A2(KEYINPUT63), .A3(new_n1228), .A4(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1224), .A2(new_n1230), .ZN(new_n1231));
  NOR3_X1   g1031(.A1(new_n1218), .A2(new_n1231), .A3(KEYINPUT61), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT62), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1216), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1234), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1233), .B1(new_n1235), .B2(new_n1214), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1227), .A2(new_n1228), .A3(new_n1229), .ZN(new_n1237));
  AOI21_X1  g1037(.A(KEYINPUT61), .B1(new_n1237), .B2(KEYINPUT62), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1224), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1194), .B1(new_n1232), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1224), .ZN(new_n1241));
  AOI21_X1  g1041(.A(KEYINPUT62), .B1(new_n1237), .B2(new_n1217), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT61), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1214), .B2(new_n1233), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1241), .B1(new_n1242), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT63), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1237), .B1(new_n1235), .B2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1243), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1245), .B(KEYINPUT126), .C1(new_n1231), .C2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1240), .A2(new_n1249), .ZN(G405));
  INV_X1    g1050(.A(G375), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1225), .B1(new_n1251), .B2(G378), .ZN(new_n1252));
  XNOR2_X1  g1052(.A(new_n1252), .B(new_n1229), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1253), .A2(KEYINPUT127), .A3(new_n1224), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT127), .B1(new_n1253), .B2(new_n1224), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n1253), .A2(new_n1224), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(G402));
endmodule


