

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U560 ( .A(KEYINPUT95), .ZN(n730) );
  XNOR2_X1 U561 ( .A(n730), .B(KEYINPUT29), .ZN(n731) );
  XNOR2_X1 U562 ( .A(n732), .B(n731), .ZN(n733) );
  NAND2_X1 U563 ( .A1(n697), .A2(n696), .ZN(n746) );
  NOR2_X1 U564 ( .A1(G651), .A2(n631), .ZN(n657) );
  XOR2_X1 U565 ( .A(KEYINPUT0), .B(G543), .Z(n631) );
  NAND2_X1 U566 ( .A1(n657), .A2(G51), .ZN(n530) );
  INV_X1 U567 ( .A(G651), .ZN(n533) );
  NOR2_X1 U568 ( .A1(G543), .A2(n533), .ZN(n527) );
  XOR2_X1 U569 ( .A(KEYINPUT66), .B(n527), .Z(n528) );
  XNOR2_X1 U570 ( .A(KEYINPUT1), .B(n528), .ZN(n652) );
  NAND2_X1 U571 ( .A1(G63), .A2(n652), .ZN(n529) );
  NAND2_X1 U572 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U573 ( .A(KEYINPUT6), .B(n531), .ZN(n539) );
  NOR2_X1 U574 ( .A1(G651), .A2(G543), .ZN(n651) );
  NAND2_X1 U575 ( .A1(n651), .A2(G89), .ZN(n532) );
  XNOR2_X1 U576 ( .A(n532), .B(KEYINPUT4), .ZN(n535) );
  NOR2_X1 U577 ( .A1(n631), .A2(n533), .ZN(n656) );
  NAND2_X1 U578 ( .A1(G76), .A2(n656), .ZN(n534) );
  NAND2_X1 U579 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U580 ( .A(KEYINPUT5), .B(n536), .ZN(n537) );
  XNOR2_X1 U581 ( .A(KEYINPUT71), .B(n537), .ZN(n538) );
  NOR2_X1 U582 ( .A1(n539), .A2(n538), .ZN(n540) );
  XOR2_X1 U583 ( .A(KEYINPUT7), .B(n540), .Z(G168) );
  XOR2_X1 U584 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U585 ( .A(G2104), .ZN(n546) );
  INV_X1 U586 ( .A(G2105), .ZN(n541) );
  NOR2_X1 U587 ( .A1(n546), .A2(n541), .ZN(n896) );
  NAND2_X1 U588 ( .A1(G113), .A2(n896), .ZN(n543) );
  NOR2_X1 U589 ( .A1(G2104), .A2(n541), .ZN(n897) );
  NAND2_X1 U590 ( .A1(G125), .A2(n897), .ZN(n542) );
  NAND2_X1 U591 ( .A1(n543), .A2(n542), .ZN(n551) );
  NOR2_X1 U592 ( .A1(G2104), .A2(G2105), .ZN(n544) );
  XOR2_X2 U593 ( .A(KEYINPUT17), .B(n544), .Z(n900) );
  NAND2_X1 U594 ( .A1(G137), .A2(n900), .ZN(n545) );
  XNOR2_X1 U595 ( .A(n545), .B(KEYINPUT64), .ZN(n549) );
  NOR2_X1 U596 ( .A1(G2105), .A2(n546), .ZN(n901) );
  NAND2_X1 U597 ( .A1(G101), .A2(n901), .ZN(n547) );
  XOR2_X1 U598 ( .A(KEYINPUT23), .B(n547), .Z(n548) );
  NAND2_X1 U599 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X2 U600 ( .A1(n551), .A2(n550), .ZN(G160) );
  NAND2_X1 U601 ( .A1(G91), .A2(n651), .ZN(n553) );
  NAND2_X1 U602 ( .A1(G78), .A2(n656), .ZN(n552) );
  NAND2_X1 U603 ( .A1(n553), .A2(n552), .ZN(n557) );
  NAND2_X1 U604 ( .A1(n657), .A2(G53), .ZN(n555) );
  NAND2_X1 U605 ( .A1(G65), .A2(n652), .ZN(n554) );
  NAND2_X1 U606 ( .A1(n555), .A2(n554), .ZN(n556) );
  OR2_X1 U607 ( .A1(n557), .A2(n556), .ZN(G299) );
  XOR2_X1 U608 ( .A(G2438), .B(G2454), .Z(n559) );
  XNOR2_X1 U609 ( .A(G2435), .B(G2430), .ZN(n558) );
  XNOR2_X1 U610 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U611 ( .A(n560), .B(KEYINPUT104), .Z(n562) );
  XNOR2_X1 U612 ( .A(G1341), .B(G1348), .ZN(n561) );
  XNOR2_X1 U613 ( .A(n562), .B(n561), .ZN(n566) );
  XOR2_X1 U614 ( .A(G2446), .B(G2451), .Z(n564) );
  XNOR2_X1 U615 ( .A(G2443), .B(G2427), .ZN(n563) );
  XNOR2_X1 U616 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U617 ( .A(n566), .B(n565), .Z(n567) );
  AND2_X1 U618 ( .A1(G14), .A2(n567), .ZN(G401) );
  NAND2_X1 U619 ( .A1(G52), .A2(n657), .ZN(n568) );
  XNOR2_X1 U620 ( .A(n568), .B(KEYINPUT67), .ZN(n575) );
  NAND2_X1 U621 ( .A1(G90), .A2(n651), .ZN(n570) );
  NAND2_X1 U622 ( .A1(G77), .A2(n656), .ZN(n569) );
  NAND2_X1 U623 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U624 ( .A(n571), .B(KEYINPUT9), .ZN(n573) );
  NAND2_X1 U625 ( .A1(G64), .A2(n652), .ZN(n572) );
  NAND2_X1 U626 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U627 ( .A1(n575), .A2(n574), .ZN(G171) );
  AND2_X1 U628 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U629 ( .A(G57), .ZN(G237) );
  NAND2_X1 U630 ( .A1(G7), .A2(G661), .ZN(n576) );
  XNOR2_X1 U631 ( .A(n576), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U632 ( .A(KEYINPUT11), .B(KEYINPUT68), .Z(n578) );
  INV_X1 U633 ( .A(G223), .ZN(n849) );
  NAND2_X1 U634 ( .A1(G567), .A2(n849), .ZN(n577) );
  XNOR2_X1 U635 ( .A(n578), .B(n577), .ZN(G234) );
  NAND2_X1 U636 ( .A1(n652), .A2(G56), .ZN(n579) );
  XOR2_X1 U637 ( .A(KEYINPUT14), .B(n579), .Z(n586) );
  NAND2_X1 U638 ( .A1(G81), .A2(n651), .ZN(n580) );
  XOR2_X1 U639 ( .A(KEYINPUT69), .B(n580), .Z(n581) );
  XNOR2_X1 U640 ( .A(n581), .B(KEYINPUT12), .ZN(n583) );
  NAND2_X1 U641 ( .A1(G68), .A2(n656), .ZN(n582) );
  NAND2_X1 U642 ( .A1(n583), .A2(n582), .ZN(n584) );
  XOR2_X1 U643 ( .A(KEYINPUT13), .B(n584), .Z(n585) );
  NOR2_X1 U644 ( .A1(n586), .A2(n585), .ZN(n588) );
  NAND2_X1 U645 ( .A1(n657), .A2(G43), .ZN(n587) );
  NAND2_X1 U646 ( .A1(n588), .A2(n587), .ZN(n952) );
  INV_X1 U647 ( .A(n952), .ZN(n708) );
  NAND2_X1 U648 ( .A1(n708), .A2(G860), .ZN(n589) );
  XNOR2_X1 U649 ( .A(KEYINPUT70), .B(n589), .ZN(G153) );
  INV_X1 U650 ( .A(G171), .ZN(G301) );
  NAND2_X1 U651 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U652 ( .A1(n657), .A2(G54), .ZN(n591) );
  NAND2_X1 U653 ( .A1(G66), .A2(n652), .ZN(n590) );
  NAND2_X1 U654 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U655 ( .A1(G92), .A2(n651), .ZN(n593) );
  NAND2_X1 U656 ( .A1(G79), .A2(n656), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U658 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U659 ( .A(n596), .B(KEYINPUT15), .ZN(n716) );
  INV_X1 U660 ( .A(G868), .ZN(n672) );
  NAND2_X1 U661 ( .A1(n716), .A2(n672), .ZN(n597) );
  NAND2_X1 U662 ( .A1(n598), .A2(n597), .ZN(G284) );
  XNOR2_X1 U663 ( .A(KEYINPUT72), .B(n672), .ZN(n599) );
  NOR2_X1 U664 ( .A1(G286), .A2(n599), .ZN(n602) );
  NOR2_X1 U665 ( .A1(G868), .A2(G299), .ZN(n600) );
  XOR2_X1 U666 ( .A(KEYINPUT73), .B(n600), .Z(n601) );
  NOR2_X1 U667 ( .A1(n602), .A2(n601), .ZN(G297) );
  INV_X1 U668 ( .A(G860), .ZN(n603) );
  NAND2_X1 U669 ( .A1(n603), .A2(G559), .ZN(n604) );
  INV_X1 U670 ( .A(n716), .ZN(n953) );
  NAND2_X1 U671 ( .A1(n604), .A2(n953), .ZN(n605) );
  XNOR2_X1 U672 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U673 ( .A1(G868), .A2(n952), .ZN(n608) );
  NAND2_X1 U674 ( .A1(n953), .A2(G868), .ZN(n606) );
  NOR2_X1 U675 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U676 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U677 ( .A1(n896), .A2(G111), .ZN(n615) );
  NAND2_X1 U678 ( .A1(G135), .A2(n900), .ZN(n610) );
  NAND2_X1 U679 ( .A1(G99), .A2(n901), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n613) );
  NAND2_X1 U681 ( .A1(n897), .A2(G123), .ZN(n611) );
  XOR2_X1 U682 ( .A(KEYINPUT18), .B(n611), .Z(n612) );
  NOR2_X1 U683 ( .A1(n613), .A2(n612), .ZN(n614) );
  NAND2_X1 U684 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U685 ( .A(KEYINPUT74), .B(n616), .Z(n1024) );
  XOR2_X1 U686 ( .A(G2096), .B(KEYINPUT75), .Z(n617) );
  XNOR2_X1 U687 ( .A(n1024), .B(n617), .ZN(n619) );
  INV_X1 U688 ( .A(G2100), .ZN(n618) );
  NAND2_X1 U689 ( .A1(n619), .A2(n618), .ZN(G156) );
  NAND2_X1 U690 ( .A1(n953), .A2(G559), .ZN(n669) );
  XNOR2_X1 U691 ( .A(n952), .B(n669), .ZN(n620) );
  NOR2_X1 U692 ( .A1(n620), .A2(G860), .ZN(n627) );
  NAND2_X1 U693 ( .A1(G93), .A2(n651), .ZN(n622) );
  NAND2_X1 U694 ( .A1(G80), .A2(n656), .ZN(n621) );
  NAND2_X1 U695 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n657), .A2(G55), .ZN(n624) );
  NAND2_X1 U697 ( .A1(G67), .A2(n652), .ZN(n623) );
  NAND2_X1 U698 ( .A1(n624), .A2(n623), .ZN(n625) );
  OR2_X1 U699 ( .A1(n626), .A2(n625), .ZN(n671) );
  XOR2_X1 U700 ( .A(n627), .B(n671), .Z(G145) );
  NAND2_X1 U701 ( .A1(G49), .A2(n657), .ZN(n629) );
  NAND2_X1 U702 ( .A1(G74), .A2(G651), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U704 ( .A(KEYINPUT76), .B(n630), .Z(n633) );
  NAND2_X1 U705 ( .A1(n631), .A2(G87), .ZN(n632) );
  NAND2_X1 U706 ( .A1(n633), .A2(n632), .ZN(n634) );
  NOR2_X1 U707 ( .A1(n634), .A2(n652), .ZN(n635) );
  XNOR2_X1 U708 ( .A(n635), .B(KEYINPUT77), .ZN(G288) );
  NAND2_X1 U709 ( .A1(G85), .A2(n651), .ZN(n637) );
  NAND2_X1 U710 ( .A1(G72), .A2(n656), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U712 ( .A(KEYINPUT65), .B(n638), .ZN(n642) );
  NAND2_X1 U713 ( .A1(n652), .A2(G60), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n657), .A2(G47), .ZN(n639) );
  AND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n641) );
  NAND2_X1 U716 ( .A1(n642), .A2(n641), .ZN(G290) );
  NAND2_X1 U717 ( .A1(G86), .A2(n651), .ZN(n644) );
  NAND2_X1 U718 ( .A1(G61), .A2(n652), .ZN(n643) );
  NAND2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U720 ( .A(KEYINPUT78), .B(n645), .ZN(n648) );
  NAND2_X1 U721 ( .A1(G73), .A2(n656), .ZN(n646) );
  XOR2_X1 U722 ( .A(KEYINPUT2), .B(n646), .Z(n647) );
  NOR2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n657), .A2(G48), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n650), .A2(n649), .ZN(G305) );
  NAND2_X1 U726 ( .A1(n651), .A2(G88), .ZN(n655) );
  NAND2_X1 U727 ( .A1(n652), .A2(G62), .ZN(n653) );
  XOR2_X1 U728 ( .A(KEYINPUT79), .B(n653), .Z(n654) );
  NAND2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n661) );
  NAND2_X1 U730 ( .A1(G75), .A2(n656), .ZN(n659) );
  NAND2_X1 U731 ( .A1(G50), .A2(n657), .ZN(n658) );
  NAND2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n660) );
  NOR2_X1 U733 ( .A1(n661), .A2(n660), .ZN(G166) );
  XNOR2_X1 U734 ( .A(G288), .B(n708), .ZN(n662) );
  XNOR2_X1 U735 ( .A(n662), .B(G290), .ZN(n665) );
  XNOR2_X1 U736 ( .A(KEYINPUT19), .B(G305), .ZN(n663) );
  XNOR2_X1 U737 ( .A(n663), .B(G299), .ZN(n664) );
  XOR2_X1 U738 ( .A(n665), .B(n664), .Z(n667) );
  XOR2_X1 U739 ( .A(G166), .B(n671), .Z(n666) );
  XNOR2_X1 U740 ( .A(n667), .B(n666), .ZN(n918) );
  XOR2_X1 U741 ( .A(n918), .B(KEYINPUT80), .Z(n668) );
  XNOR2_X1 U742 ( .A(n669), .B(n668), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n670), .A2(G868), .ZN(n674) );
  NAND2_X1 U744 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U745 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U747 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U748 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U750 ( .A1(n678), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U752 ( .A1(G69), .A2(G120), .ZN(n679) );
  NOR2_X1 U753 ( .A1(G237), .A2(n679), .ZN(n680) );
  NAND2_X1 U754 ( .A1(G108), .A2(n680), .ZN(n854) );
  NAND2_X1 U755 ( .A1(G567), .A2(n854), .ZN(n687) );
  XOR2_X1 U756 ( .A(KEYINPUT22), .B(KEYINPUT81), .Z(n682) );
  NAND2_X1 U757 ( .A1(G132), .A2(G82), .ZN(n681) );
  XNOR2_X1 U758 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U759 ( .A1(n683), .A2(G218), .ZN(n684) );
  XNOR2_X1 U760 ( .A(KEYINPUT82), .B(n684), .ZN(n685) );
  NAND2_X1 U761 ( .A1(n685), .A2(G96), .ZN(n853) );
  NAND2_X1 U762 ( .A1(G2106), .A2(n853), .ZN(n686) );
  NAND2_X1 U763 ( .A1(n687), .A2(n686), .ZN(n855) );
  NAND2_X1 U764 ( .A1(G661), .A2(G483), .ZN(n688) );
  NOR2_X1 U765 ( .A1(n855), .A2(n688), .ZN(n852) );
  NAND2_X1 U766 ( .A1(n852), .A2(G36), .ZN(G176) );
  NAND2_X1 U767 ( .A1(G138), .A2(n900), .ZN(n690) );
  NAND2_X1 U768 ( .A1(G102), .A2(n901), .ZN(n689) );
  NAND2_X1 U769 ( .A1(n690), .A2(n689), .ZN(n694) );
  NAND2_X1 U770 ( .A1(G114), .A2(n896), .ZN(n692) );
  NAND2_X1 U771 ( .A1(G126), .A2(n897), .ZN(n691) );
  NAND2_X1 U772 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U773 ( .A1(n694), .A2(n693), .ZN(G164) );
  XNOR2_X1 U774 ( .A(KEYINPUT83), .B(G166), .ZN(G303) );
  XNOR2_X1 U775 ( .A(G1986), .B(G290), .ZN(n957) );
  NOR2_X1 U776 ( .A1(G164), .A2(G1384), .ZN(n697) );
  NAND2_X1 U777 ( .A1(G160), .A2(G40), .ZN(n695) );
  NOR2_X1 U778 ( .A1(n697), .A2(n695), .ZN(n843) );
  NAND2_X1 U779 ( .A1(n957), .A2(n843), .ZN(n830) );
  XOR2_X1 U780 ( .A(G1981), .B(G305), .Z(n960) );
  XOR2_X1 U781 ( .A(G1961), .B(KEYINPUT90), .Z(n985) );
  INV_X1 U782 ( .A(n695), .ZN(n696) );
  NAND2_X1 U783 ( .A1(n985), .A2(n746), .ZN(n699) );
  INV_X1 U784 ( .A(n746), .ZN(n719) );
  XNOR2_X1 U785 ( .A(G2078), .B(KEYINPUT25), .ZN(n934) );
  NAND2_X1 U786 ( .A1(n719), .A2(n934), .ZN(n698) );
  NAND2_X1 U787 ( .A1(n699), .A2(n698), .ZN(n739) );
  AND2_X1 U788 ( .A1(n739), .A2(G171), .ZN(n700) );
  XNOR2_X1 U789 ( .A(KEYINPUT91), .B(n700), .ZN(n734) );
  XNOR2_X1 U790 ( .A(G1996), .B(KEYINPUT92), .ZN(n940) );
  NAND2_X1 U791 ( .A1(n719), .A2(n940), .ZN(n701) );
  XNOR2_X1 U792 ( .A(n701), .B(KEYINPUT26), .ZN(n703) );
  AND2_X1 U793 ( .A1(n746), .A2(G1341), .ZN(n702) );
  NAND2_X1 U794 ( .A1(KEYINPUT26), .A2(n702), .ZN(n706) );
  NAND2_X1 U795 ( .A1(n703), .A2(n706), .ZN(n705) );
  INV_X1 U796 ( .A(KEYINPUT93), .ZN(n704) );
  NAND2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n710) );
  NAND2_X1 U798 ( .A1(n706), .A2(KEYINPUT93), .ZN(n707) );
  AND2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n709) );
  AND2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n714) );
  NAND2_X1 U801 ( .A1(G1348), .A2(n746), .ZN(n712) );
  NAND2_X1 U802 ( .A1(G2067), .A2(n719), .ZN(n711) );
  NAND2_X1 U803 ( .A1(n712), .A2(n711), .ZN(n715) );
  NOR2_X1 U804 ( .A1(n716), .A2(n715), .ZN(n713) );
  NOR2_X1 U805 ( .A1(n714), .A2(n713), .ZN(n718) );
  AND2_X1 U806 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U807 ( .A1(n718), .A2(n717), .ZN(n724) );
  NAND2_X1 U808 ( .A1(n719), .A2(G2072), .ZN(n720) );
  XOR2_X1 U809 ( .A(KEYINPUT27), .B(n720), .Z(n722) );
  NAND2_X1 U810 ( .A1(G1956), .A2(n746), .ZN(n721) );
  NAND2_X1 U811 ( .A1(n722), .A2(n721), .ZN(n726) );
  NOR2_X1 U812 ( .A1(G299), .A2(n726), .ZN(n723) );
  NOR2_X1 U813 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U814 ( .A(KEYINPUT94), .B(n725), .ZN(n729) );
  NAND2_X1 U815 ( .A1(G299), .A2(n726), .ZN(n727) );
  XOR2_X1 U816 ( .A(n727), .B(KEYINPUT28), .Z(n728) );
  NOR2_X1 U817 ( .A1(n729), .A2(n728), .ZN(n732) );
  NAND2_X1 U818 ( .A1(n734), .A2(n733), .ZN(n744) );
  NAND2_X1 U819 ( .A1(G8), .A2(n746), .ZN(n792) );
  NOR2_X1 U820 ( .A1(G1966), .A2(n792), .ZN(n760) );
  NOR2_X1 U821 ( .A1(n746), .A2(G2084), .ZN(n735) );
  XNOR2_X1 U822 ( .A(n735), .B(KEYINPUT89), .ZN(n756) );
  NAND2_X1 U823 ( .A1(G8), .A2(n756), .ZN(n736) );
  NOR2_X1 U824 ( .A1(n760), .A2(n736), .ZN(n737) );
  XOR2_X1 U825 ( .A(KEYINPUT30), .B(n737), .Z(n738) );
  NOR2_X1 U826 ( .A1(G168), .A2(n738), .ZN(n741) );
  NOR2_X1 U827 ( .A1(G171), .A2(n739), .ZN(n740) );
  NOR2_X1 U828 ( .A1(n741), .A2(n740), .ZN(n742) );
  XOR2_X1 U829 ( .A(KEYINPUT31), .B(n742), .Z(n743) );
  NAND2_X1 U830 ( .A1(n744), .A2(n743), .ZN(n758) );
  NAND2_X1 U831 ( .A1(n758), .A2(G286), .ZN(n745) );
  XNOR2_X1 U832 ( .A(n745), .B(KEYINPUT96), .ZN(n753) );
  NOR2_X1 U833 ( .A1(G2090), .A2(n746), .ZN(n748) );
  NOR2_X1 U834 ( .A1(G1971), .A2(n792), .ZN(n747) );
  NOR2_X1 U835 ( .A1(n748), .A2(n747), .ZN(n749) );
  XOR2_X1 U836 ( .A(KEYINPUT97), .B(n749), .Z(n750) );
  NAND2_X1 U837 ( .A1(n750), .A2(G303), .ZN(n751) );
  XNOR2_X1 U838 ( .A(KEYINPUT98), .B(n751), .ZN(n752) );
  NAND2_X1 U839 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U840 ( .A1(n754), .A2(G8), .ZN(n755) );
  XNOR2_X1 U841 ( .A(KEYINPUT32), .B(n755), .ZN(n783) );
  INV_X1 U842 ( .A(n756), .ZN(n757) );
  NAND2_X1 U843 ( .A1(G8), .A2(n757), .ZN(n762) );
  INV_X1 U844 ( .A(n758), .ZN(n759) );
  NOR2_X1 U845 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n762), .A2(n761), .ZN(n784) );
  AND2_X1 U847 ( .A1(G288), .A2(G1976), .ZN(n966) );
  NOR2_X1 U848 ( .A1(n966), .A2(n792), .ZN(n772) );
  AND2_X1 U849 ( .A1(n784), .A2(n772), .ZN(n764) );
  INV_X1 U850 ( .A(KEYINPUT99), .ZN(n763) );
  AND2_X1 U851 ( .A1(n764), .A2(n763), .ZN(n770) );
  NOR2_X1 U852 ( .A1(G1976), .A2(G288), .ZN(n774) );
  NAND2_X1 U853 ( .A1(n774), .A2(KEYINPUT33), .ZN(n765) );
  NAND2_X1 U854 ( .A1(n763), .A2(n765), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n774), .A2(KEYINPUT99), .ZN(n766) );
  NAND2_X1 U856 ( .A1(n767), .A2(n766), .ZN(n768) );
  NOR2_X1 U857 ( .A1(n792), .A2(n768), .ZN(n779) );
  INV_X1 U858 ( .A(n779), .ZN(n769) );
  AND2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n783), .A2(n771), .ZN(n781) );
  INV_X1 U861 ( .A(n772), .ZN(n775) );
  NOR2_X1 U862 ( .A1(G1971), .A2(G303), .ZN(n773) );
  NOR2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n972) );
  OR2_X1 U864 ( .A1(n775), .A2(n972), .ZN(n776) );
  NOR2_X1 U865 ( .A1(KEYINPUT99), .A2(n776), .ZN(n777) );
  NOR2_X1 U866 ( .A1(n777), .A2(KEYINPUT33), .ZN(n778) );
  OR2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  AND2_X1 U869 ( .A1(n960), .A2(n782), .ZN(n797) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n788) );
  NOR2_X1 U871 ( .A1(G2090), .A2(G303), .ZN(n785) );
  NAND2_X1 U872 ( .A1(G8), .A2(n785), .ZN(n786) );
  XNOR2_X1 U873 ( .A(n786), .B(KEYINPUT100), .ZN(n787) );
  NAND2_X1 U874 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U875 ( .A1(n789), .A2(n792), .ZN(n795) );
  NOR2_X1 U876 ( .A1(G1981), .A2(G305), .ZN(n790) );
  XOR2_X1 U877 ( .A(n790), .B(KEYINPUT24), .Z(n791) );
  NOR2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U879 ( .A(n793), .B(KEYINPUT88), .Z(n794) );
  NAND2_X1 U880 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U881 ( .A1(n797), .A2(n796), .ZN(n828) );
  NAND2_X1 U882 ( .A1(G105), .A2(n901), .ZN(n798) );
  XNOR2_X1 U883 ( .A(n798), .B(KEYINPUT86), .ZN(n799) );
  XNOR2_X1 U884 ( .A(n799), .B(KEYINPUT38), .ZN(n801) );
  NAND2_X1 U885 ( .A1(G141), .A2(n900), .ZN(n800) );
  NAND2_X1 U886 ( .A1(n801), .A2(n800), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G129), .A2(n897), .ZN(n802) );
  XNOR2_X1 U888 ( .A(KEYINPUT85), .B(n802), .ZN(n803) );
  NOR2_X1 U889 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U890 ( .A1(n896), .A2(G117), .ZN(n805) );
  NAND2_X1 U891 ( .A1(n806), .A2(n805), .ZN(n910) );
  AND2_X1 U892 ( .A1(n910), .A2(G1996), .ZN(n814) );
  INV_X1 U893 ( .A(G1991), .ZN(n831) );
  NAND2_X1 U894 ( .A1(G131), .A2(n900), .ZN(n808) );
  NAND2_X1 U895 ( .A1(G95), .A2(n901), .ZN(n807) );
  NAND2_X1 U896 ( .A1(n808), .A2(n807), .ZN(n812) );
  NAND2_X1 U897 ( .A1(G107), .A2(n896), .ZN(n810) );
  NAND2_X1 U898 ( .A1(G119), .A2(n897), .ZN(n809) );
  NAND2_X1 U899 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U900 ( .A1(n812), .A2(n811), .ZN(n895) );
  NOR2_X1 U901 ( .A1(n831), .A2(n895), .ZN(n813) );
  NOR2_X1 U902 ( .A1(n814), .A2(n813), .ZN(n1029) );
  XNOR2_X1 U903 ( .A(KEYINPUT87), .B(n843), .ZN(n815) );
  NOR2_X1 U904 ( .A1(n1029), .A2(n815), .ZN(n834) );
  INV_X1 U905 ( .A(n834), .ZN(n826) );
  XNOR2_X1 U906 ( .A(KEYINPUT37), .B(G2067), .ZN(n840) );
  NAND2_X1 U907 ( .A1(G140), .A2(n900), .ZN(n817) );
  NAND2_X1 U908 ( .A1(G104), .A2(n901), .ZN(n816) );
  NAND2_X1 U909 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U910 ( .A(KEYINPUT34), .B(n818), .ZN(n824) );
  NAND2_X1 U911 ( .A1(n897), .A2(G128), .ZN(n819) );
  XNOR2_X1 U912 ( .A(n819), .B(KEYINPUT84), .ZN(n821) );
  NAND2_X1 U913 ( .A1(G116), .A2(n896), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n821), .A2(n820), .ZN(n822) );
  XOR2_X1 U915 ( .A(KEYINPUT35), .B(n822), .Z(n823) );
  NOR2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U917 ( .A(KEYINPUT36), .B(n825), .ZN(n915) );
  NOR2_X1 U918 ( .A1(n840), .A2(n915), .ZN(n1022) );
  NAND2_X1 U919 ( .A1(n843), .A2(n1022), .ZN(n838) );
  NAND2_X1 U920 ( .A1(n826), .A2(n838), .ZN(n827) );
  NOR2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n847) );
  NOR2_X1 U923 ( .A1(G1996), .A2(n910), .ZN(n1015) );
  NOR2_X1 U924 ( .A1(G1986), .A2(G290), .ZN(n832) );
  AND2_X1 U925 ( .A1(n831), .A2(n895), .ZN(n1023) );
  NOR2_X1 U926 ( .A1(n832), .A2(n1023), .ZN(n833) );
  NOR2_X1 U927 ( .A1(n834), .A2(n833), .ZN(n835) );
  NOR2_X1 U928 ( .A1(n1015), .A2(n835), .ZN(n836) );
  XOR2_X1 U929 ( .A(n836), .B(KEYINPUT101), .Z(n837) );
  XNOR2_X1 U930 ( .A(n837), .B(KEYINPUT39), .ZN(n839) );
  NAND2_X1 U931 ( .A1(n839), .A2(n838), .ZN(n841) );
  NAND2_X1 U932 ( .A1(n840), .A2(n915), .ZN(n1019) );
  NAND2_X1 U933 ( .A1(n841), .A2(n1019), .ZN(n842) );
  XNOR2_X1 U934 ( .A(KEYINPUT102), .B(n842), .ZN(n844) );
  NAND2_X1 U935 ( .A1(n844), .A2(n843), .ZN(n845) );
  XOR2_X1 U936 ( .A(KEYINPUT103), .B(n845), .Z(n846) );
  NAND2_X1 U937 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U938 ( .A(KEYINPUT40), .B(n848), .ZN(G329) );
  NAND2_X1 U939 ( .A1(G2106), .A2(n849), .ZN(G217) );
  AND2_X1 U940 ( .A1(G15), .A2(G2), .ZN(n850) );
  NAND2_X1 U941 ( .A1(G661), .A2(n850), .ZN(G259) );
  NAND2_X1 U942 ( .A1(G3), .A2(G1), .ZN(n851) );
  NAND2_X1 U943 ( .A1(n852), .A2(n851), .ZN(G188) );
  INV_X1 U945 ( .A(G132), .ZN(G219) );
  INV_X1 U946 ( .A(G120), .ZN(G236) );
  INV_X1 U947 ( .A(G96), .ZN(G221) );
  INV_X1 U948 ( .A(G82), .ZN(G220) );
  INV_X1 U949 ( .A(G69), .ZN(G235) );
  NOR2_X1 U950 ( .A1(n854), .A2(n853), .ZN(G325) );
  INV_X1 U951 ( .A(G325), .ZN(G261) );
  INV_X1 U952 ( .A(n855), .ZN(G319) );
  XOR2_X1 U953 ( .A(G2100), .B(KEYINPUT106), .Z(n857) );
  XNOR2_X1 U954 ( .A(KEYINPUT105), .B(KEYINPUT43), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U956 ( .A(KEYINPUT42), .B(G2090), .Z(n859) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2072), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U959 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U960 ( .A(G2678), .B(G2096), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n865) );
  XOR2_X1 U962 ( .A(G2078), .B(G2084), .Z(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(G227) );
  XOR2_X1 U964 ( .A(G1986), .B(G1961), .Z(n867) );
  XNOR2_X1 U965 ( .A(G1981), .B(G1966), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U967 ( .A(G1971), .B(G1976), .Z(n869) );
  XNOR2_X1 U968 ( .A(G1991), .B(G1996), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U970 ( .A(n871), .B(n870), .Z(n873) );
  XNOR2_X1 U971 ( .A(G2474), .B(KEYINPUT41), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(n875) );
  XOR2_X1 U973 ( .A(G1956), .B(KEYINPUT107), .Z(n874) );
  XNOR2_X1 U974 ( .A(n875), .B(n874), .ZN(G229) );
  NAND2_X1 U975 ( .A1(G124), .A2(n897), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n876), .B(KEYINPUT44), .ZN(n879) );
  NAND2_X1 U977 ( .A1(G100), .A2(n901), .ZN(n877) );
  XNOR2_X1 U978 ( .A(n877), .B(KEYINPUT108), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n883) );
  NAND2_X1 U980 ( .A1(G136), .A2(n900), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G112), .A2(n896), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U983 ( .A1(n883), .A2(n882), .ZN(G162) );
  XOR2_X1 U984 ( .A(KEYINPUT110), .B(KEYINPUT46), .Z(n893) );
  NAND2_X1 U985 ( .A1(G115), .A2(n896), .ZN(n885) );
  NAND2_X1 U986 ( .A1(G127), .A2(n897), .ZN(n884) );
  NAND2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n886) );
  XNOR2_X1 U988 ( .A(n886), .B(KEYINPUT47), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G103), .A2(n901), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n891) );
  NAND2_X1 U991 ( .A1(G139), .A2(n900), .ZN(n889) );
  XNOR2_X1 U992 ( .A(KEYINPUT109), .B(n889), .ZN(n890) );
  NOR2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n1008) );
  XNOR2_X1 U994 ( .A(n1008), .B(KEYINPUT48), .ZN(n892) );
  XNOR2_X1 U995 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U996 ( .A(n895), .B(n894), .ZN(n914) );
  XNOR2_X1 U997 ( .A(G160), .B(G162), .ZN(n908) );
  NAND2_X1 U998 ( .A1(G118), .A2(n896), .ZN(n899) );
  NAND2_X1 U999 ( .A1(G130), .A2(n897), .ZN(n898) );
  NAND2_X1 U1000 ( .A1(n899), .A2(n898), .ZN(n906) );
  NAND2_X1 U1001 ( .A1(G142), .A2(n900), .ZN(n903) );
  NAND2_X1 U1002 ( .A1(G106), .A2(n901), .ZN(n902) );
  NAND2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1004 ( .A(KEYINPUT45), .B(n904), .Z(n905) );
  NOR2_X1 U1005 ( .A1(n906), .A2(n905), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n1024), .B(n909), .ZN(n912) );
  XOR2_X1 U1008 ( .A(n910), .B(G164), .Z(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n914), .B(n913), .ZN(n916) );
  XOR2_X1 U1011 ( .A(n916), .B(n915), .Z(n917) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n917), .ZN(G395) );
  XNOR2_X1 U1013 ( .A(G171), .B(G286), .ZN(n919) );
  XNOR2_X1 U1014 ( .A(n919), .B(n918), .ZN(n920) );
  XNOR2_X1 U1015 ( .A(n920), .B(n953), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n921), .ZN(G397) );
  NOR2_X1 U1017 ( .A1(G227), .A2(G229), .ZN(n922) );
  XOR2_X1 U1018 ( .A(KEYINPUT49), .B(n922), .Z(n923) );
  NAND2_X1 U1019 ( .A1(G319), .A2(n923), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(G401), .A2(n924), .ZN(n927) );
  NOR2_X1 U1021 ( .A1(G395), .A2(G397), .ZN(n925) );
  XOR2_X1 U1022 ( .A(KEYINPUT111), .B(n925), .Z(n926) );
  NAND2_X1 U1023 ( .A1(n927), .A2(n926), .ZN(G225) );
  INV_X1 U1024 ( .A(G225), .ZN(G308) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1026 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n1041) );
  XNOR2_X1 U1027 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n928) );
  XNOR2_X1 U1028 ( .A(n928), .B(G34), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(G2084), .B(n929), .ZN(n947) );
  XNOR2_X1 U1030 ( .A(G2090), .B(G35), .ZN(n945) );
  XNOR2_X1 U1031 ( .A(G25), .B(G1991), .ZN(n930) );
  XNOR2_X1 U1032 ( .A(n930), .B(KEYINPUT117), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(G2067), .B(G26), .ZN(n932) );
  XNOR2_X1 U1034 ( .A(G33), .B(G2072), .ZN(n931) );
  NOR2_X1 U1035 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1036 ( .A1(G28), .A2(n933), .ZN(n937) );
  XOR2_X1 U1037 ( .A(G27), .B(n934), .Z(n935) );
  XNOR2_X1 U1038 ( .A(KEYINPUT118), .B(n935), .ZN(n936) );
  NOR2_X1 U1039 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1040 ( .A1(n939), .A2(n938), .ZN(n942) );
  XNOR2_X1 U1041 ( .A(G32), .B(n940), .ZN(n941) );
  NOR2_X1 U1042 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1043 ( .A(KEYINPUT53), .B(n943), .ZN(n944) );
  NOR2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(n948), .B(KEYINPUT120), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(n949), .B(KEYINPUT55), .ZN(n950) );
  NOR2_X1 U1048 ( .A1(G29), .A2(n950), .ZN(n1005) );
  XNOR2_X1 U1049 ( .A(G16), .B(KEYINPUT56), .ZN(n974) );
  INV_X1 U1050 ( .A(G1341), .ZN(n951) );
  XNOR2_X1 U1051 ( .A(n952), .B(n951), .ZN(n959) );
  XNOR2_X1 U1052 ( .A(G1348), .B(n953), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(G1971), .A2(G303), .ZN(n954) );
  NAND2_X1 U1054 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n970) );
  XNOR2_X1 U1057 ( .A(G1966), .B(G168), .ZN(n961) );
  NAND2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(n962), .B(KEYINPUT57), .ZN(n968) );
  XOR2_X1 U1060 ( .A(G299), .B(G1956), .Z(n964) );
  XNOR2_X1 U1061 ( .A(G171), .B(G1961), .ZN(n963) );
  NAND2_X1 U1062 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1063 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1065 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n1003) );
  INV_X1 U1068 ( .A(G16), .ZN(n1001) );
  XNOR2_X1 U1069 ( .A(G1348), .B(KEYINPUT59), .ZN(n975) );
  XNOR2_X1 U1070 ( .A(n975), .B(G4), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(G1981), .B(G6), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(G1956), .B(G20), .ZN(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n982) );
  XOR2_X1 U1075 ( .A(KEYINPUT121), .B(G1341), .Z(n980) );
  XNOR2_X1 U1076 ( .A(G19), .B(n980), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(KEYINPUT122), .B(n983), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(n984), .B(KEYINPUT60), .ZN(n996) );
  XOR2_X1 U1080 ( .A(n985), .B(G5), .Z(n994) );
  XNOR2_X1 U1081 ( .A(KEYINPUT123), .B(G1971), .ZN(n986) );
  XNOR2_X1 U1082 ( .A(n986), .B(G22), .ZN(n991) );
  XNOR2_X1 U1083 ( .A(G1986), .B(KEYINPUT124), .ZN(n987) );
  XNOR2_X1 U1084 ( .A(n987), .B(G24), .ZN(n989) );
  XNOR2_X1 U1085 ( .A(G23), .B(G1976), .ZN(n988) );
  NOR2_X1 U1086 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1087 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1088 ( .A(n992), .B(KEYINPUT58), .ZN(n993) );
  NOR2_X1 U1089 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1090 ( .A1(n996), .A2(n995), .ZN(n998) );
  XNOR2_X1 U1091 ( .A(G21), .B(G1966), .ZN(n997) );
  NOR2_X1 U1092 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1093 ( .A(KEYINPUT61), .B(n999), .ZN(n1000) );
  NAND2_X1 U1094 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1095 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(G11), .A2(n1006), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(n1007), .B(KEYINPUT125), .ZN(n1039) );
  XNOR2_X1 U1099 ( .A(G2072), .B(n1008), .ZN(n1011) );
  XNOR2_X1 U1100 ( .A(G164), .B(G2078), .ZN(n1009) );
  XNOR2_X1 U1101 ( .A(n1009), .B(KEYINPUT116), .ZN(n1010) );
  NAND2_X1 U1102 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XNOR2_X1 U1103 ( .A(n1012), .B(KEYINPUT50), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(G2090), .B(G162), .ZN(n1013) );
  XNOR2_X1 U1105 ( .A(n1013), .B(KEYINPUT115), .ZN(n1014) );
  NOR2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1107 ( .A(KEYINPUT51), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  NAND2_X1 U1109 ( .A1(n1020), .A2(n1019), .ZN(n1033) );
  XOR2_X1 U1110 ( .A(G160), .B(G2084), .Z(n1021) );
  NOR2_X1 U1111 ( .A1(n1022), .A2(n1021), .ZN(n1027) );
  NOR2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1113 ( .A(n1025), .B(KEYINPUT112), .ZN(n1026) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1115 ( .A(KEYINPUT113), .B(n1028), .ZN(n1030) );
  NAND2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XNOR2_X1 U1117 ( .A(KEYINPUT114), .B(n1031), .ZN(n1032) );
  NOR2_X1 U1118 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1119 ( .A(KEYINPUT52), .B(n1034), .ZN(n1036) );
  INV_X1 U1120 ( .A(KEYINPUT55), .ZN(n1035) );
  NAND2_X1 U1121 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1122 ( .A1(n1037), .A2(G29), .ZN(n1038) );
  NAND2_X1 U1123 ( .A1(n1039), .A2(n1038), .ZN(n1040) );
  XNOR2_X1 U1124 ( .A(n1041), .B(n1040), .ZN(G150) );
  INV_X1 U1125 ( .A(G150), .ZN(G311) );
endmodule

