//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 1 0 1 0 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n800, new_n801, new_n802, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1052, new_n1053, new_n1054;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(G169gat), .B(G197gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT95), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT17), .ZN(new_n209));
  INV_X1    g008(.A(G36gat), .ZN(new_n210));
  AND2_X1   g009(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT15), .ZN(new_n214));
  INV_X1    g013(.A(G29gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n215), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n214), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT94), .ZN(new_n218));
  INV_X1    g017(.A(G43gat), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n218), .B1(new_n219), .B2(G50gat), .ZN(new_n220));
  AOI22_X1  g019(.A1(new_n213), .A2(new_n216), .B1(new_n214), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G43gat), .B(G50gat), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n217), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n220), .A2(new_n214), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT14), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n215), .ZN(new_n226));
  NAND2_X1  g025(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n227));
  AOI21_X1  g026(.A(G36gat), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n215), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n224), .B(new_n222), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  OAI211_X1 g030(.A(new_n208), .B(new_n209), .C1(new_n223), .C2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n224), .B1(new_n228), .B2(new_n229), .ZN(new_n233));
  INV_X1    g032(.A(new_n222), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n226), .A2(new_n227), .ZN(new_n235));
  AOI21_X1  g034(.A(new_n229), .B1(new_n235), .B2(new_n210), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n233), .A2(new_n234), .B1(new_n236), .B2(new_n214), .ZN(new_n237));
  NAND2_X1  g036(.A1(KEYINPUT95), .A2(KEYINPUT17), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n208), .A2(new_n209), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n237), .A2(new_n230), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n232), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G15gat), .B(G22gat), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n242), .A2(G1gat), .ZN(new_n243));
  AOI21_X1  g042(.A(G8gat), .B1(new_n243), .B2(KEYINPUT96), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT16), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n242), .B1(new_n245), .B2(G1gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n243), .B(new_n246), .C1(KEYINPUT96), .C2(G8gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n241), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(G229gat), .A2(G233gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n230), .ZN(new_n253));
  INV_X1    g052(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(new_n249), .A3(new_n248), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n251), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT18), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n250), .A2(new_n253), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n252), .B(KEYINPUT13), .Z(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n251), .A2(KEYINPUT18), .A3(new_n255), .A4(new_n252), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n207), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n258), .A2(new_n264), .A3(new_n262), .A4(new_n207), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(G169gat), .A2(G176gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(KEYINPUT23), .ZN(new_n270));
  NAND2_X1  g069(.A1(G169gat), .A2(G176gat), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OR2_X1    g071(.A1(new_n269), .A2(KEYINPUT23), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n275), .A2(KEYINPUT66), .ZN(new_n276));
  INV_X1    g075(.A(G183gat), .ZN(new_n277));
  INV_X1    g076(.A(G190gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT66), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n279), .B(new_n280), .C1(new_n274), .C2(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(new_n272), .B(new_n273), .C1(new_n276), .C2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(KEYINPUT65), .B(KEYINPUT25), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT67), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n270), .A2(new_n287), .A3(new_n271), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n270), .B2(new_n271), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g089(.A(KEYINPUT25), .B1(new_n269), .B2(KEYINPUT23), .ZN(new_n291));
  AND2_X1   g090(.A1(new_n279), .A2(new_n280), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(new_n275), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n286), .A2(new_n294), .ZN(new_n295));
  OR2_X1    g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT26), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n296), .A2(new_n297), .A3(new_n271), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n269), .A2(KEYINPUT26), .ZN(new_n299));
  NAND2_X1  g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT28), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n277), .A2(KEYINPUT27), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(KEYINPUT68), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(new_n278), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT27), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G183gat), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT68), .B1(new_n303), .B2(new_n307), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n302), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n303), .A2(new_n307), .ZN(new_n310));
  INV_X1    g109(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(KEYINPUT28), .A3(new_n278), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n301), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT69), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI211_X1 g114(.A(KEYINPUT69), .B(new_n301), .C1(new_n309), .C2(new_n312), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n295), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OR2_X1    g116(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(KEYINPUT70), .A2(G127gat), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n318), .A2(KEYINPUT71), .A3(G134gat), .A4(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n321));
  INV_X1    g120(.A(G113gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(G120gat), .ZN(new_n323));
  INV_X1    g122(.A(G120gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(G113gat), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n321), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n318), .A2(G134gat), .A3(new_n319), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT71), .ZN(new_n328));
  INV_X1    g127(.A(G127gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n328), .B1(new_n329), .B2(G134gat), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n320), .B(new_n326), .C1(new_n327), .C2(new_n330), .ZN(new_n331));
  XOR2_X1   g130(.A(G127gat), .B(G134gat), .Z(new_n332));
  OR2_X1    g131(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT72), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(new_n333), .A3(KEYINPUT72), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n317), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n337), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT72), .B1(new_n331), .B2(new_n333), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n301), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT68), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n310), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g144(.A(G190gat), .B1(new_n303), .B2(KEYINPUT68), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT28), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n310), .A2(new_n302), .A3(G190gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n343), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(KEYINPUT69), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n313), .A2(new_n314), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n342), .A2(new_n352), .A3(new_n295), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n339), .A2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(G227gat), .ZN(new_n355));
  INV_X1    g154(.A(G233gat), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(KEYINPUT64), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT32), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT33), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(G15gat), .B(G43gat), .Z(new_n363));
  XNOR2_X1  g162(.A(G71gat), .B(G99gat), .ZN(new_n364));
  XNOR2_X1  g163(.A(new_n363), .B(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n360), .A2(new_n362), .A3(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n358), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n367), .B1(new_n339), .B2(new_n353), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n365), .B1(new_n368), .B2(KEYINPUT33), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT32), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g171(.A(new_n339), .B(new_n353), .C1(new_n355), .C2(new_n356), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT34), .ZN(new_n374));
  AND2_X1   g173(.A1(new_n339), .A2(new_n353), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n358), .A2(KEYINPUT34), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n374), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n366), .A2(KEYINPUT73), .A3(new_n372), .A4(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n369), .A2(new_n371), .ZN(new_n380));
  AOI221_X4 g179(.A(new_n370), .B1(KEYINPUT33), .B2(new_n365), .C1(new_n354), .C2(new_n358), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT73), .ZN(new_n382));
  AOI22_X1  g181(.A1(KEYINPUT34), .A2(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n383));
  OAI22_X1  g182(.A1(new_n380), .A2(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT36), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n383), .B1(new_n380), .B2(new_n381), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n366), .A2(new_n372), .A3(new_n378), .ZN(new_n388));
  XOR2_X1   g187(.A(KEYINPUT74), .B(KEYINPUT36), .Z(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n386), .A2(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G8gat), .B(G36gat), .ZN(new_n392));
  XNOR2_X1  g191(.A(G64gat), .B(G92gat), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n392), .B(new_n393), .Z(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  AND2_X1   g194(.A1(G211gat), .A2(G218gat), .ZN(new_n396));
  NOR2_X1   g195(.A1(G211gat), .A2(G218gat), .ZN(new_n397));
  OAI21_X1  g196(.A(KEYINPUT76), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(G211gat), .ZN(new_n399));
  INV_X1    g198(.A(G218gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT76), .ZN(new_n402));
  NAND2_X1  g201(.A1(G211gat), .A2(G218gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  OR2_X1    g204(.A1(G197gat), .A2(G204gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(G197gat), .A2(G204gat), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT22), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n406), .A2(new_n407), .B1(new_n408), .B2(new_n403), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n405), .A2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT77), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT77), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n405), .A2(new_n412), .A3(new_n409), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT75), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n405), .B1(new_n414), .B2(new_n409), .ZN(new_n415));
  OR2_X1    g214(.A1(new_n409), .A2(new_n414), .ZN(new_n416));
  AOI22_X1  g215(.A1(new_n411), .A2(new_n413), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AND2_X1   g216(.A1(G226gat), .A2(G233gat), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n295), .A2(new_n418), .A3(new_n349), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n283), .A2(new_n285), .B1(new_n290), .B2(new_n293), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n420), .B1(new_n350), .B2(new_n351), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n418), .A2(KEYINPUT29), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n417), .B(new_n419), .C1(new_n421), .C2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n352), .A2(new_n418), .A3(new_n295), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n295), .A2(new_n349), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(new_n422), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n417), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n395), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  AOI22_X1  g229(.A1(new_n421), .A2(new_n418), .B1(new_n427), .B2(new_n422), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n424), .B(new_n394), .C1(new_n431), .C2(new_n417), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(KEYINPUT30), .A3(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n425), .A2(new_n429), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT30), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n394), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT6), .ZN(new_n438));
  XNOR2_X1  g237(.A(G155gat), .B(G162gat), .ZN(new_n439));
  XOR2_X1   g238(.A(G141gat), .B(G148gat), .Z(new_n440));
  XOR2_X1   g239(.A(KEYINPUT78), .B(KEYINPUT2), .Z(new_n441));
  AOI21_X1  g240(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n439), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT2), .ZN(new_n444));
  XNOR2_X1  g243(.A(KEYINPUT79), .B(G162gat), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n444), .B1(new_n445), .B2(G155gat), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT80), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  AND2_X1   g246(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n448));
  NOR2_X1   g247(.A1(KEYINPUT79), .A2(G162gat), .ZN(new_n449));
  OAI21_X1  g248(.A(G155gat), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT2), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT80), .ZN(new_n452));
  NAND4_X1  g251(.A1(new_n451), .A2(new_n452), .A3(new_n439), .A4(new_n440), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n442), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n334), .ZN(new_n455));
  AND3_X1   g254(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT4), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT4), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n336), .A2(new_n454), .A3(new_n337), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n456), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(G225gat), .A2(G233gat), .ZN(new_n460));
  XOR2_X1   g259(.A(new_n460), .B(KEYINPUT81), .Z(new_n461));
  NAND2_X1  g260(.A1(new_n447), .A2(new_n453), .ZN(new_n462));
  INV_X1    g261(.A(new_n442), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n455), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n454), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n461), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT5), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n459), .A2(new_n468), .A3(KEYINPUT83), .A4(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT83), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n458), .A2(new_n457), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT4), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n461), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n334), .B1(new_n454), .B2(new_n466), .ZN(new_n476));
  AOI211_X1 g275(.A(KEYINPUT3), .B(new_n442), .C1(new_n447), .C2(new_n453), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n469), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n471), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n470), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n458), .A2(KEYINPUT4), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(KEYINPUT82), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT82), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n458), .A2(new_n484), .A3(KEYINPUT4), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n468), .A3(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n454), .B(new_n455), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n469), .B1(new_n487), .B2(new_n461), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n480), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G1gat), .B(G29gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(KEYINPUT0), .ZN(new_n492));
  XNOR2_X1  g291(.A(G57gat), .B(G85gat), .ZN(new_n493));
  XOR2_X1   g292(.A(new_n492), .B(new_n493), .Z(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT84), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n470), .A2(new_n479), .B1(new_n486), .B2(new_n488), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n497), .B1(new_n498), .B2(new_n494), .ZN(new_n499));
  AND4_X1   g298(.A1(new_n497), .A2(new_n480), .A3(new_n494), .A4(new_n489), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n438), .B(new_n496), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(new_n496), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n437), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G78gat), .B(G106gat), .ZN(new_n505));
  INV_X1    g304(.A(G50gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n505), .B(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT29), .B1(new_n454), .B2(new_n466), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n411), .A2(new_n413), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n415), .A2(new_n416), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT86), .B1(new_n508), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT29), .B1(new_n509), .B2(new_n510), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n464), .B1(new_n513), .B2(KEYINPUT3), .ZN(new_n514));
  INV_X1    g313(.A(G228gat), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(new_n356), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT86), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n517), .B(new_n417), .C1(new_n477), .C2(KEYINPUT29), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n512), .A2(new_n514), .A3(new_n516), .A4(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n405), .A2(new_n412), .A3(new_n409), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n412), .B1(new_n405), .B2(new_n409), .ZN(new_n521));
  OAI22_X1  g320(.A1(new_n520), .A2(new_n521), .B1(new_n405), .B2(new_n409), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT29), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n454), .B1(new_n524), .B2(new_n466), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n511), .B1(new_n467), .B2(new_n523), .ZN(new_n526));
  OAI22_X1  g325(.A1(new_n525), .A2(new_n526), .B1(new_n515), .B2(new_n356), .ZN(new_n527));
  INV_X1    g326(.A(G22gat), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n519), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n528), .B1(new_n519), .B2(new_n527), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n507), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n519), .A2(new_n527), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n532), .A2(G22gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n519), .A2(new_n527), .A3(new_n528), .ZN(new_n534));
  INV_X1    g333(.A(new_n507), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n531), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n531), .B2(new_n536), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n391), .B1(new_n504), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT87), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT87), .ZN(new_n544));
  OAI211_X1 g343(.A(new_n544), .B(new_n391), .C1(new_n504), .C2(new_n541), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT84), .B1(new_n490), .B2(new_n495), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n498), .A2(new_n497), .A3(new_n494), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT6), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT88), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n498), .B2(new_n494), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n490), .A2(KEYINPUT88), .A3(new_n495), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g351(.A1(new_n548), .A2(new_n552), .B1(KEYINPUT6), .B2(new_n502), .ZN(new_n553));
  XOR2_X1   g352(.A(KEYINPUT90), .B(KEYINPUT37), .Z(new_n554));
  AOI21_X1  g353(.A(new_n394), .B1(new_n434), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT38), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n511), .B(new_n419), .C1(new_n421), .C2(new_n423), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n557), .B(KEYINPUT37), .C1(new_n431), .C2(new_n511), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n555), .A2(new_n556), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n559), .A2(new_n432), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT37), .B1(new_n425), .B2(new_n429), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n556), .B1(new_n555), .B2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n553), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n565), .A2(new_n334), .A3(new_n467), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n566), .A2(new_n472), .A3(new_n473), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT39), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n461), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n475), .B1(new_n459), .B2(new_n566), .ZN(new_n570));
  OAI21_X1  g369(.A(KEYINPUT39), .B1(new_n487), .B2(new_n461), .ZN(new_n571));
  OAI211_X1 g370(.A(new_n569), .B(new_n494), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT40), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n437), .A2(new_n550), .A3(new_n551), .A4(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(KEYINPUT89), .B1(new_n572), .B2(new_n573), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n495), .B1(new_n570), .B2(new_n568), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT89), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n567), .A2(new_n461), .ZN(new_n579));
  INV_X1    g378(.A(new_n571), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT40), .A4(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(new_n576), .A2(new_n582), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n575), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n564), .A2(new_n541), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n543), .A2(new_n545), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n385), .B1(new_n538), .B2(new_n539), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT92), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT92), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n385), .B(new_n589), .C1(new_n538), .C2(new_n539), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n588), .A2(new_n504), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT35), .ZN(new_n592));
  AND3_X1   g391(.A1(new_n387), .A2(new_n388), .A3(KEYINPUT91), .ZN(new_n593));
  AOI21_X1  g392(.A(KEYINPUT91), .B1(new_n387), .B2(new_n388), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n437), .A2(KEYINPUT35), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(new_n538), .B2(new_n539), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n553), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n592), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n268), .B1(new_n586), .B2(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n501), .A2(new_n503), .ZN(new_n603));
  XOR2_X1   g402(.A(G190gat), .B(G218gat), .Z(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G99gat), .B(G106gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  OR2_X1    g406(.A1(KEYINPUT100), .A2(G92gat), .ZN(new_n608));
  INV_X1    g407(.A(G85gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(KEYINPUT100), .A2(G92gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G99gat), .A2(G106gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT8), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G85gat), .A2(G92gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(KEYINPUT99), .A2(KEYINPUT7), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n607), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT101), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n615), .A2(KEYINPUT99), .A3(KEYINPUT7), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n616), .A2(G85gat), .A3(G92gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n622), .A2(new_n606), .A3(new_n611), .A4(new_n613), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n618), .A2(new_n619), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n622), .A2(new_n611), .A3(new_n613), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(KEYINPUT101), .A3(new_n607), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n624), .A2(KEYINPUT102), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(KEYINPUT102), .B1(new_n624), .B2(new_n626), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n241), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT103), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n241), .B(KEYINPUT103), .C1(new_n627), .C2(new_n628), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n623), .A2(new_n619), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT8), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n636), .B1(G99gat), .B2(G106gat), .ZN(new_n637));
  AND2_X1   g436(.A1(KEYINPUT100), .A2(G92gat), .ZN(new_n638));
  NOR2_X1   g437(.A1(KEYINPUT100), .A2(G92gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n637), .B1(new_n640), .B2(new_n609), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n606), .B1(new_n641), .B2(new_n622), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n635), .A2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n626), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n634), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n624), .A2(KEYINPUT102), .A3(new_n626), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n254), .A3(new_n646), .ZN(new_n647));
  AND2_X1   g446(.A1(G232gat), .A2(G233gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT41), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n605), .B1(new_n633), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n648), .A2(KEYINPUT41), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT98), .ZN(new_n655));
  XNOR2_X1  g454(.A(G134gat), .B(G162gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n633), .A2(new_n605), .A3(new_n651), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n653), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n657), .ZN(new_n660));
  AOI211_X1 g459(.A(new_n604), .B(new_n650), .C1(new_n631), .C2(new_n632), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n660), .B1(new_n661), .B2(new_n652), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(G64gat), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n664), .A2(G57gat), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(G57gat), .ZN(new_n666));
  INV_X1    g465(.A(G71gat), .ZN(new_n667));
  INV_X1    g466(.A(G78gat), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI22_X1  g468(.A1(new_n665), .A2(new_n666), .B1(new_n669), .B2(KEYINPUT9), .ZN(new_n670));
  XOR2_X1   g469(.A(G71gat), .B(G78gat), .Z(new_n671));
  XNOR2_X1  g470(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT21), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(G127gat), .B(G155gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n250), .B1(new_n673), .B2(new_n672), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(G231gat), .A2(G233gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT97), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(G183gat), .B(G211gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n678), .B(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n663), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(G120gat), .B(G148gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(G176gat), .B(G204gat), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n688), .B(new_n689), .Z(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(G230gat), .A2(G233gat), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT10), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n672), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n645), .A2(new_n646), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n624), .A2(new_n672), .A3(new_n626), .ZN(new_n697));
  INV_X1    g496(.A(new_n671), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n670), .B(new_n698), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(new_n618), .A3(new_n623), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n697), .A2(new_n700), .A3(new_n694), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n693), .B1(new_n696), .B2(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(KEYINPUT105), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704));
  AOI211_X1 g503(.A(new_n704), .B(new_n693), .C1(new_n696), .C2(new_n701), .ZN(new_n705));
  NOR2_X1   g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n697), .A2(new_n700), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(new_n693), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n691), .B1(new_n706), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n701), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n711), .B1(new_n712), .B2(new_n692), .ZN(new_n713));
  AOI211_X1 g512(.A(KEYINPUT104), .B(new_n693), .C1(new_n696), .C2(new_n701), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n709), .A2(new_n691), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n687), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n602), .A2(new_n603), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g522(.A1(new_n602), .A2(new_n721), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n437), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n725), .A2(G8gat), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT16), .B(G8gat), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n725), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT42), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n729), .B1(KEYINPUT42), .B2(new_n728), .ZN(G1325gat));
  INV_X1    g529(.A(G15gat), .ZN(new_n731));
  INV_X1    g530(.A(new_n595), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n724), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n391), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n724), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n733), .B1(new_n735), .B2(new_n731), .ZN(G1326gat));
  NAND2_X1  g535(.A1(new_n724), .A2(new_n540), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT43), .B(G22gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n737), .B(new_n738), .ZN(G1327gat));
  INV_X1    g538(.A(new_n663), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n740), .A2(new_n685), .A3(new_n718), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n602), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n742), .A2(new_n215), .A3(new_n603), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n743), .B(KEYINPUT45), .ZN(new_n744));
  OAI22_X1  g543(.A1(new_n575), .A2(new_n583), .B1(new_n538), .B2(new_n539), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n745), .B1(new_n553), .B2(new_n563), .ZN(new_n746));
  OR2_X1    g545(.A1(new_n746), .A2(new_n542), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT107), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n601), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n591), .A2(KEYINPUT35), .B1(new_n598), .B2(new_n599), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n746), .A2(new_n542), .ZN(new_n751));
  OAI21_X1  g550(.A(KEYINPUT107), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n740), .A2(KEYINPUT44), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n749), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n740), .B1(new_n586), .B2(new_n601), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  XOR2_X1   g556(.A(new_n685), .B(KEYINPUT106), .Z(new_n758));
  INV_X1    g557(.A(new_n268), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n758), .A2(new_n759), .A3(new_n719), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n761), .A2(new_n603), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n744), .B1(new_n762), .B2(new_n215), .ZN(G1328gat));
  NAND3_X1  g562(.A1(new_n742), .A2(new_n210), .A3(new_n437), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(KEYINPUT46), .Z(new_n765));
  AND2_X1   g564(.A1(new_n761), .A2(new_n437), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n765), .B1(new_n766), .B2(new_n210), .ZN(G1329gat));
  NAND3_X1  g566(.A1(new_n742), .A2(new_n219), .A3(new_n732), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(new_n770));
  AND3_X1   g569(.A1(new_n757), .A2(new_n734), .A3(new_n760), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n770), .B(KEYINPUT47), .C1(new_n771), .C2(new_n219), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT47), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n768), .B(KEYINPUT108), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n771), .A2(new_n219), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n772), .A2(new_n776), .ZN(G1330gat));
  NAND3_X1  g576(.A1(new_n742), .A2(new_n506), .A3(new_n540), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n757), .A2(new_n540), .A3(new_n760), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n779), .B2(new_n506), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT109), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT48), .B1(new_n778), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n780), .B(new_n782), .ZN(G1331gat));
  AND2_X1   g582(.A1(new_n749), .A2(new_n752), .ZN(new_n784));
  NOR4_X1   g583(.A1(new_n759), .A2(new_n663), .A3(new_n719), .A4(new_n686), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n603), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g587(.A1(new_n784), .A2(new_n785), .ZN(new_n789));
  INV_X1    g588(.A(new_n437), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n791), .A2(new_n664), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  OR3_X1    g593(.A1(new_n789), .A2(KEYINPUT110), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT110), .B1(new_n789), .B2(new_n794), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n791), .A2(new_n664), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n797), .B(new_n798), .ZN(G1333gat));
  NAND3_X1  g598(.A1(new_n786), .A2(new_n667), .A3(new_n732), .ZN(new_n800));
  OAI21_X1  g599(.A(G71gat), .B1(new_n789), .B2(new_n391), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XOR2_X1   g601(.A(new_n802), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g602(.A1(new_n789), .A2(new_n541), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(new_n668), .ZN(G1335gat));
  INV_X1    g604(.A(KEYINPUT111), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n268), .A2(new_n686), .ZN(new_n807));
  NOR2_X1   g606(.A1(new_n807), .A2(new_n719), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n757), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n806), .B1(new_n757), .B2(new_n808), .ZN(new_n811));
  INV_X1    g610(.A(new_n603), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n740), .A2(new_n807), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n814), .B1(new_n750), .B2(new_n751), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT51), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g616(.A(KEYINPUT51), .B(new_n814), .C1(new_n750), .C2(new_n751), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n603), .A2(new_n609), .A3(new_n718), .ZN(new_n821));
  XOR2_X1   g620(.A(new_n821), .B(KEYINPUT112), .Z(new_n822));
  OAI22_X1  g621(.A1(new_n813), .A2(new_n609), .B1(new_n820), .B2(new_n822), .ZN(G1336gat));
  NAND2_X1  g622(.A1(new_n819), .A2(new_n718), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n824), .A2(G92gat), .A3(new_n790), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(KEYINPUT52), .ZN(new_n826));
  INV_X1    g625(.A(new_n640), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n749), .A2(new_n752), .A3(new_n753), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n586), .A2(new_n601), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n755), .B1(new_n829), .B2(new_n663), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n808), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n827), .B1(new_n831), .B2(new_n790), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n826), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n831), .A2(KEYINPUT111), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n437), .A3(new_n809), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n825), .B1(new_n835), .B2(new_n827), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(G1337gat));
  NOR3_X1   g637(.A1(new_n810), .A2(new_n811), .A3(new_n391), .ZN(new_n839));
  XNOR2_X1  g638(.A(KEYINPUT113), .B(G99gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n732), .A2(new_n840), .ZN(new_n841));
  OAI22_X1  g640(.A1(new_n839), .A2(new_n840), .B1(new_n824), .B2(new_n841), .ZN(G1338gat));
  NOR2_X1   g641(.A1(new_n541), .A2(G106gat), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n819), .A2(new_n718), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT114), .ZN(new_n845));
  AOI21_X1  g644(.A(KEYINPUT53), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n819), .A2(KEYINPUT114), .A3(new_n718), .A4(new_n843), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n831), .B2(new_n541), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n757), .A2(KEYINPUT115), .A3(new_n540), .A4(new_n808), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(G106gat), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n848), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(new_n844), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n834), .A2(new_n540), .A3(new_n809), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n854), .B1(new_n855), .B2(G106gat), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT53), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(G1339gat));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n690), .B1(new_n706), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n696), .A2(new_n693), .A3(new_n701), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n861), .A2(KEYINPUT54), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT116), .B1(new_n715), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n699), .A2(KEYINPUT10), .ZN(new_n864));
  NOR3_X1   g663(.A1(new_n627), .A2(new_n628), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g664(.A1(new_n697), .A2(new_n700), .A3(new_n694), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n692), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(KEYINPUT104), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n702), .A2(new_n711), .ZN(new_n869));
  AND4_X1   g668(.A1(KEYINPUT116), .A2(new_n868), .A3(new_n862), .A4(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n860), .B1(new_n863), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n268), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(KEYINPUT55), .B(new_n860), .C1(new_n863), .C2(new_n870), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n874), .A2(KEYINPUT117), .A3(new_n717), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT117), .B1(new_n874), .B2(new_n717), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n250), .A2(new_n253), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n878), .B1(new_n250), .B2(new_n241), .ZN(new_n879));
  OAI22_X1  g678(.A1(new_n879), .A2(new_n252), .B1(new_n260), .B2(new_n261), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n206), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n266), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n882), .B1(new_n710), .B2(new_n717), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n663), .B1(new_n877), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n266), .A2(KEYINPUT118), .A3(new_n881), .ZN(new_n888));
  AND4_X1   g687(.A1(new_n659), .A2(new_n887), .A3(new_n662), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n871), .A2(new_n872), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n717), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n874), .A2(KEYINPUT117), .A3(new_n717), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n758), .B1(new_n885), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n720), .A2(new_n759), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n588), .A2(new_n590), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n900), .A2(new_n603), .A3(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(new_n437), .ZN(new_n903));
  AOI21_X1  g702(.A(G113gat), .B1(new_n903), .B2(new_n759), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n595), .A2(new_n540), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n900), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n603), .A2(new_n790), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n268), .A2(new_n322), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n904), .B1(new_n908), .B2(new_n909), .ZN(G1340gat));
  AOI21_X1  g709(.A(G120gat), .B1(new_n903), .B2(new_n718), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n719), .A2(new_n324), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n911), .B1(new_n908), .B2(new_n912), .ZN(G1341gat));
  NAND2_X1  g712(.A1(new_n318), .A2(new_n319), .ZN(new_n914));
  INV_X1    g713(.A(new_n908), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n915), .B2(new_n758), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n903), .A2(new_n318), .A3(new_n319), .A4(new_n685), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1342gat));
  OAI21_X1  g717(.A(G134gat), .B1(new_n915), .B2(new_n740), .ZN(new_n919));
  OR3_X1    g718(.A1(new_n740), .A2(G134gat), .A3(new_n437), .ZN(new_n920));
  OR3_X1    g719(.A1(new_n902), .A2(KEYINPUT56), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g720(.A(KEYINPUT56), .B1(new_n902), .B2(new_n920), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(G1343gat));
  NOR2_X1   g722(.A1(new_n907), .A2(new_n734), .ZN(new_n924));
  AOI21_X1  g723(.A(KEYINPUT57), .B1(new_n900), .B2(new_n540), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n868), .A2(new_n862), .A3(new_n869), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT116), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n715), .A2(KEYINPUT116), .A3(new_n862), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT55), .B1(new_n930), .B2(new_n860), .ZN(new_n931));
  NAND4_X1  g730(.A1(new_n659), .A2(new_n887), .A3(new_n662), .A4(new_n888), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n933), .B1(new_n875), .B2(new_n876), .ZN(new_n934));
  INV_X1    g733(.A(new_n717), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n867), .A2(new_n704), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n702), .A2(KEYINPUT105), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n936), .A2(new_n859), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n691), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n939), .B1(new_n928), .B2(new_n929), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n935), .B1(new_n940), .B2(KEYINPUT55), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n883), .B1(new_n941), .B2(new_n873), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n934), .B1(new_n663), .B2(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n898), .B1(new_n943), .B2(new_n686), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT57), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n944), .A2(new_n945), .A3(new_n541), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n924), .B1(new_n925), .B2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(new_n759), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G141gat), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n391), .A2(new_n540), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n951), .A2(new_n437), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n900), .A2(new_n603), .A3(new_n952), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n268), .A2(G141gat), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  XNOR2_X1  g755(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n950), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(KEYINPUT119), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT119), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n954), .A2(new_n960), .A3(new_n955), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n962), .B1(G141gat), .B2(new_n949), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT58), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n958), .B1(new_n963), .B2(new_n964), .ZN(G1344gat));
  OR3_X1    g764(.A1(new_n953), .A2(G148gat), .A3(new_n719), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT59), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n941), .A2(new_n873), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n663), .B1(new_n969), .B2(new_n884), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n968), .B1(new_n970), .B2(new_n896), .ZN(new_n971));
  OAI211_X1 g770(.A(new_n934), .B(KEYINPUT121), .C1(new_n663), .C2(new_n942), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n971), .A2(new_n686), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n973), .A2(new_n899), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n541), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n685), .B1(new_n943), .B2(new_n968), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n898), .B1(new_n977), .B2(new_n972), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(KEYINPUT122), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT57), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n541), .A2(new_n945), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n900), .A2(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(new_n982), .ZN(new_n983));
  OAI211_X1 g782(.A(new_n718), .B(new_n924), .C1(new_n980), .C2(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n967), .B1(new_n984), .B2(G148gat), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n967), .A2(G148gat), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n986), .B1(new_n948), .B2(new_n718), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n966), .B1(new_n985), .B2(new_n987), .ZN(G1345gat));
  INV_X1    g787(.A(G155gat), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n947), .A2(new_n989), .A3(new_n758), .ZN(new_n990));
  OAI21_X1  g789(.A(KEYINPUT123), .B1(new_n953), .B2(new_n686), .ZN(new_n991));
  NOR3_X1   g790(.A1(new_n953), .A2(KEYINPUT123), .A3(new_n686), .ZN(new_n992));
  NOR2_X1   g791(.A1(new_n992), .A2(G155gat), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n990), .B1(new_n991), .B2(new_n993), .ZN(G1346gat));
  OAI21_X1  g793(.A(new_n445), .B1(new_n947), .B2(new_n740), .ZN(new_n995));
  OR2_X1    g794(.A1(new_n740), .A2(new_n445), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n995), .B1(new_n953), .B2(new_n996), .ZN(G1347gat));
  NOR2_X1   g796(.A1(new_n603), .A2(new_n790), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n900), .A2(new_n905), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g798(.A(G169gat), .B1(new_n999), .B2(new_n268), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT124), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n603), .B1(new_n897), .B2(new_n899), .ZN(new_n1002));
  AND2_X1   g801(.A1(new_n901), .A2(new_n437), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g803(.A(new_n1004), .ZN(new_n1005));
  NOR2_X1   g804(.A1(new_n268), .A2(G169gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1001), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NOR4_X1   g806(.A1(new_n1004), .A2(KEYINPUT124), .A3(G169gat), .A4(new_n268), .ZN(new_n1008));
  OAI21_X1  g807(.A(new_n1000), .B1(new_n1007), .B2(new_n1008), .ZN(G1348gat));
  OAI21_X1  g808(.A(G176gat), .B1(new_n999), .B2(new_n719), .ZN(new_n1010));
  OR2_X1    g809(.A1(new_n719), .A2(G176gat), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1010), .B1(new_n1004), .B2(new_n1011), .ZN(G1349gat));
  NOR2_X1   g811(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n1005), .A2(new_n311), .A3(new_n685), .ZN(new_n1014));
  OAI21_X1  g813(.A(G183gat), .B1(new_n999), .B2(new_n758), .ZN(new_n1015));
  AOI21_X1  g814(.A(new_n1013), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g815(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n1017));
  XOR2_X1   g816(.A(new_n1016), .B(new_n1017), .Z(G1350gat));
  OAI21_X1  g817(.A(G190gat), .B1(new_n999), .B2(new_n740), .ZN(new_n1019));
  INV_X1    g818(.A(KEYINPUT126), .ZN(new_n1020));
  AND2_X1   g819(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g820(.A(KEYINPUT61), .ZN(new_n1022));
  NOR2_X1   g821(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g822(.A(new_n1023), .B1(new_n1020), .B2(new_n1019), .ZN(new_n1024));
  NOR3_X1   g823(.A1(new_n1004), .A2(G190gat), .A3(new_n740), .ZN(new_n1025));
  AOI21_X1  g824(.A(new_n1025), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1026));
  NAND2_X1  g825(.A1(new_n1024), .A2(new_n1026), .ZN(G1351gat));
  AND4_X1   g826(.A1(new_n437), .A2(new_n1002), .A3(new_n540), .A4(new_n391), .ZN(new_n1028));
  AOI21_X1  g827(.A(G197gat), .B1(new_n1028), .B2(new_n759), .ZN(new_n1029));
  OAI21_X1  g828(.A(new_n540), .B1(new_n978), .B2(KEYINPUT122), .ZN(new_n1030));
  NOR2_X1   g829(.A1(new_n974), .A2(new_n975), .ZN(new_n1031));
  OAI21_X1  g830(.A(new_n945), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1032), .A2(new_n982), .ZN(new_n1033));
  NOR3_X1   g832(.A1(new_n734), .A2(new_n603), .A3(new_n790), .ZN(new_n1034));
  AND2_X1   g833(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AND2_X1   g834(.A1(new_n759), .A2(G197gat), .ZN(new_n1036));
  AOI21_X1  g835(.A(new_n1029), .B1(new_n1035), .B2(new_n1036), .ZN(G1352gat));
  OAI211_X1 g836(.A(new_n718), .B(new_n1034), .C1(new_n980), .C2(new_n983), .ZN(new_n1038));
  NAND2_X1  g837(.A1(new_n1038), .A2(KEYINPUT127), .ZN(new_n1039));
  INV_X1    g838(.A(KEYINPUT127), .ZN(new_n1040));
  NAND4_X1  g839(.A1(new_n1033), .A2(new_n1040), .A3(new_n718), .A4(new_n1034), .ZN(new_n1041));
  NAND3_X1  g840(.A1(new_n1039), .A2(G204gat), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g841(.A(G204gat), .ZN(new_n1043));
  NAND3_X1  g842(.A1(new_n1028), .A2(new_n1043), .A3(new_n718), .ZN(new_n1044));
  XOR2_X1   g843(.A(new_n1044), .B(KEYINPUT62), .Z(new_n1045));
  NAND2_X1  g844(.A1(new_n1042), .A2(new_n1045), .ZN(G1353gat));
  NAND3_X1  g845(.A1(new_n1028), .A2(new_n399), .A3(new_n685), .ZN(new_n1047));
  OAI211_X1 g846(.A(new_n685), .B(new_n1034), .C1(new_n980), .C2(new_n983), .ZN(new_n1048));
  AND3_X1   g847(.A1(new_n1048), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1049));
  AOI21_X1  g848(.A(KEYINPUT63), .B1(new_n1048), .B2(G211gat), .ZN(new_n1050));
  OAI21_X1  g849(.A(new_n1047), .B1(new_n1049), .B2(new_n1050), .ZN(G1354gat));
  NAND3_X1  g850(.A1(new_n1033), .A2(new_n663), .A3(new_n1034), .ZN(new_n1052));
  NAND2_X1  g851(.A1(new_n1052), .A2(G218gat), .ZN(new_n1053));
  NAND3_X1  g852(.A1(new_n1028), .A2(new_n400), .A3(new_n663), .ZN(new_n1054));
  NAND2_X1  g853(.A1(new_n1053), .A2(new_n1054), .ZN(G1355gat));
endmodule


