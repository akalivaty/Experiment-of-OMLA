

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U557 ( .A1(n549), .A2(n548), .ZN(n550) );
  OR2_X1 U558 ( .A1(n822), .A2(n525), .ZN(n524) );
  AND2_X1 U559 ( .A1(n954), .A2(n836), .ZN(n525) );
  XOR2_X1 U560 ( .A(KEYINPUT103), .B(n782), .Z(n526) );
  XNOR2_X1 U561 ( .A(KEYINPUT31), .B(KEYINPUT99), .ZN(n740) );
  XNOR2_X1 U562 ( .A(n741), .B(n740), .ZN(n742) );
  INV_X1 U563 ( .A(n729), .ZN(n744) );
  NOR2_X1 U564 ( .A1(G651), .A2(n661), .ZN(n656) );
  OR2_X1 U565 ( .A1(n823), .A2(n524), .ZN(n839) );
  XOR2_X1 U566 ( .A(KEYINPUT15), .B(n604), .Z(n952) );
  XNOR2_X1 U567 ( .A(KEYINPUT85), .B(n550), .ZN(G164) );
  NOR2_X1 U568 ( .A1(G543), .A2(G651), .ZN(n527) );
  XNOR2_X1 U569 ( .A(n527), .B(KEYINPUT64), .ZN(n649) );
  NAND2_X1 U570 ( .A1(G89), .A2(n649), .ZN(n528) );
  XNOR2_X1 U571 ( .A(n528), .B(KEYINPUT4), .ZN(n530) );
  XOR2_X1 U572 ( .A(KEYINPUT0), .B(G543), .Z(n661) );
  INV_X1 U573 ( .A(G651), .ZN(n532) );
  NOR2_X2 U574 ( .A1(n661), .A2(n532), .ZN(n648) );
  NAND2_X1 U575 ( .A1(G76), .A2(n648), .ZN(n529) );
  NAND2_X1 U576 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U577 ( .A(n531), .B(KEYINPUT5), .ZN(n539) );
  NOR2_X1 U578 ( .A1(G543), .A2(n532), .ZN(n534) );
  XNOR2_X1 U579 ( .A(KEYINPUT1), .B(KEYINPUT67), .ZN(n533) );
  XNOR2_X1 U580 ( .A(n534), .B(n533), .ZN(n660) );
  NAND2_X1 U581 ( .A1(G63), .A2(n660), .ZN(n536) );
  NAND2_X1 U582 ( .A1(G51), .A2(n656), .ZN(n535) );
  NAND2_X1 U583 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U584 ( .A(KEYINPUT6), .B(n537), .Z(n538) );
  NAND2_X1 U585 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U586 ( .A(n540), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U587 ( .A(G168), .B(KEYINPUT8), .Z(n541) );
  XNOR2_X1 U588 ( .A(KEYINPUT74), .B(n541), .ZN(G286) );
  INV_X1 U589 ( .A(G2104), .ZN(n545) );
  AND2_X1 U590 ( .A1(n545), .A2(G2105), .ZN(n873) );
  NAND2_X1 U591 ( .A1(G126), .A2(n873), .ZN(n544) );
  OR2_X1 U592 ( .A1(G2104), .A2(G2105), .ZN(n542) );
  XNOR2_X2 U593 ( .A(KEYINPUT17), .B(n542), .ZN(n869) );
  NAND2_X1 U594 ( .A1(G138), .A2(n869), .ZN(n543) );
  NAND2_X1 U595 ( .A1(n544), .A2(n543), .ZN(n549) );
  AND2_X1 U596 ( .A1(G2104), .A2(G2105), .ZN(n874) );
  NAND2_X1 U597 ( .A1(G114), .A2(n874), .ZN(n547) );
  NOR2_X1 U598 ( .A1(G2105), .A2(n545), .ZN(n870) );
  NAND2_X1 U599 ( .A1(G102), .A2(n870), .ZN(n546) );
  NAND2_X1 U600 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U601 ( .A(G2427), .B(G2435), .Z(n552) );
  XNOR2_X1 U602 ( .A(G2454), .B(G2443), .ZN(n551) );
  XNOR2_X1 U603 ( .A(n552), .B(n551), .ZN(n559) );
  XOR2_X1 U604 ( .A(G2451), .B(KEYINPUT107), .Z(n554) );
  XNOR2_X1 U605 ( .A(G2430), .B(G2438), .ZN(n553) );
  XNOR2_X1 U606 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U607 ( .A(n555), .B(G2446), .Z(n557) );
  XNOR2_X1 U608 ( .A(G1341), .B(G1348), .ZN(n556) );
  XNOR2_X1 U609 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U610 ( .A(n559), .B(n558), .ZN(n560) );
  AND2_X1 U611 ( .A1(n560), .A2(G14), .ZN(G401) );
  AND2_X1 U612 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U613 ( .A1(G111), .A2(n874), .ZN(n562) );
  NAND2_X1 U614 ( .A1(G99), .A2(n870), .ZN(n561) );
  NAND2_X1 U615 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U616 ( .A1(G123), .A2(n873), .ZN(n563) );
  XNOR2_X1 U617 ( .A(n563), .B(KEYINPUT77), .ZN(n564) );
  XNOR2_X1 U618 ( .A(n564), .B(KEYINPUT18), .ZN(n565) );
  NOR2_X1 U619 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U620 ( .A1(n869), .A2(G135), .ZN(n567) );
  NAND2_X1 U621 ( .A1(n568), .A2(n567), .ZN(n1011) );
  XNOR2_X1 U622 ( .A(G2096), .B(n1011), .ZN(n569) );
  OR2_X1 U623 ( .A1(G2100), .A2(n569), .ZN(G156) );
  INV_X1 U624 ( .A(G57), .ZN(G237) );
  INV_X1 U625 ( .A(G132), .ZN(G219) );
  NAND2_X1 U626 ( .A1(G64), .A2(n660), .ZN(n571) );
  NAND2_X1 U627 ( .A1(G52), .A2(n656), .ZN(n570) );
  NAND2_X1 U628 ( .A1(n571), .A2(n570), .ZN(n577) );
  NAND2_X1 U629 ( .A1(n648), .A2(G77), .ZN(n573) );
  NAND2_X1 U630 ( .A1(G90), .A2(n649), .ZN(n572) );
  NAND2_X1 U631 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U632 ( .A(KEYINPUT9), .B(n574), .Z(n575) );
  XNOR2_X1 U633 ( .A(KEYINPUT68), .B(n575), .ZN(n576) );
  NOR2_X1 U634 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U635 ( .A(KEYINPUT69), .B(n578), .Z(G171) );
  INV_X1 U636 ( .A(G171), .ZN(G301) );
  NAND2_X1 U637 ( .A1(G137), .A2(n869), .ZN(n579) );
  XOR2_X1 U638 ( .A(KEYINPUT65), .B(n579), .Z(n582) );
  NAND2_X1 U639 ( .A1(G101), .A2(n870), .ZN(n580) );
  XOR2_X1 U640 ( .A(KEYINPUT23), .B(n580), .Z(n581) );
  NAND2_X1 U641 ( .A1(n582), .A2(n581), .ZN(n694) );
  NAND2_X1 U642 ( .A1(G125), .A2(n873), .ZN(n584) );
  NAND2_X1 U643 ( .A1(G113), .A2(n874), .ZN(n583) );
  NAND2_X1 U644 ( .A1(n584), .A2(n583), .ZN(n692) );
  NOR2_X1 U645 ( .A1(n694), .A2(n692), .ZN(G160) );
  NAND2_X1 U646 ( .A1(G7), .A2(G661), .ZN(n585) );
  XNOR2_X1 U647 ( .A(n585), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U648 ( .A(G223), .ZN(n841) );
  NAND2_X1 U649 ( .A1(n841), .A2(G567), .ZN(n586) );
  XOR2_X1 U650 ( .A(KEYINPUT11), .B(n586), .Z(G234) );
  NAND2_X1 U651 ( .A1(n660), .A2(G56), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(KEYINPUT14), .ZN(n589) );
  NAND2_X1 U653 ( .A1(G43), .A2(n656), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n596) );
  NAND2_X1 U655 ( .A1(G81), .A2(n649), .ZN(n590) );
  XNOR2_X1 U656 ( .A(n590), .B(KEYINPUT12), .ZN(n592) );
  NAND2_X1 U657 ( .A1(G68), .A2(n648), .ZN(n591) );
  NAND2_X1 U658 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U659 ( .A(KEYINPUT13), .B(n593), .Z(n594) );
  XNOR2_X1 U660 ( .A(KEYINPUT72), .B(n594), .ZN(n595) );
  NOR2_X2 U661 ( .A1(n596), .A2(n595), .ZN(n951) );
  NAND2_X1 U662 ( .A1(n951), .A2(G860), .ZN(G153) );
  NAND2_X1 U663 ( .A1(G868), .A2(G301), .ZN(n606) );
  NAND2_X1 U664 ( .A1(G92), .A2(n649), .ZN(n603) );
  NAND2_X1 U665 ( .A1(G66), .A2(n660), .ZN(n598) );
  NAND2_X1 U666 ( .A1(G54), .A2(n656), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G79), .A2(n648), .ZN(n599) );
  XNOR2_X1 U669 ( .A(KEYINPUT73), .B(n599), .ZN(n600) );
  NOR2_X1 U670 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n603), .A2(n602), .ZN(n604) );
  INV_X1 U672 ( .A(G868), .ZN(n620) );
  NAND2_X1 U673 ( .A1(n952), .A2(n620), .ZN(n605) );
  NAND2_X1 U674 ( .A1(n606), .A2(n605), .ZN(G284) );
  NAND2_X1 U675 ( .A1(G65), .A2(n660), .ZN(n608) );
  NAND2_X1 U676 ( .A1(G53), .A2(n656), .ZN(n607) );
  NAND2_X1 U677 ( .A1(n608), .A2(n607), .ZN(n612) );
  NAND2_X1 U678 ( .A1(n648), .A2(G78), .ZN(n610) );
  NAND2_X1 U679 ( .A1(G91), .A2(n649), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n610), .A2(n609), .ZN(n611) );
  NOR2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n955) );
  XOR2_X1 U682 ( .A(n955), .B(KEYINPUT70), .Z(G299) );
  NAND2_X1 U683 ( .A1(G868), .A2(G286), .ZN(n614) );
  NAND2_X1 U684 ( .A1(G299), .A2(n620), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n614), .A2(n613), .ZN(G297) );
  INV_X1 U686 ( .A(G860), .ZN(n624) );
  NAND2_X1 U687 ( .A1(G559), .A2(n624), .ZN(n615) );
  XOR2_X1 U688 ( .A(KEYINPUT75), .B(n615), .Z(n616) );
  INV_X1 U689 ( .A(n952), .ZN(n697) );
  NAND2_X1 U690 ( .A1(n616), .A2(n697), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n617), .B(KEYINPUT16), .ZN(n618) );
  XNOR2_X1 U692 ( .A(KEYINPUT76), .B(n618), .ZN(G148) );
  NAND2_X1 U693 ( .A1(n697), .A2(G868), .ZN(n619) );
  NOR2_X1 U694 ( .A1(G559), .A2(n619), .ZN(n622) );
  AND2_X1 U695 ( .A1(n620), .A2(n951), .ZN(n621) );
  NOR2_X1 U696 ( .A1(n622), .A2(n621), .ZN(G282) );
  NAND2_X1 U697 ( .A1(G559), .A2(n697), .ZN(n623) );
  XNOR2_X1 U698 ( .A(n623), .B(n951), .ZN(n672) );
  NAND2_X1 U699 ( .A1(n624), .A2(n672), .ZN(n632) );
  NAND2_X1 U700 ( .A1(n648), .A2(G80), .ZN(n625) );
  XNOR2_X1 U701 ( .A(n625), .B(KEYINPUT78), .ZN(n627) );
  NAND2_X1 U702 ( .A1(G67), .A2(n660), .ZN(n626) );
  NAND2_X1 U703 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U704 ( .A1(n656), .A2(G55), .ZN(n629) );
  NAND2_X1 U705 ( .A1(G93), .A2(n649), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U707 ( .A1(n631), .A2(n630), .ZN(n674) );
  XOR2_X1 U708 ( .A(n632), .B(n674), .Z(G145) );
  NAND2_X1 U709 ( .A1(n648), .A2(G72), .ZN(n634) );
  NAND2_X1 U710 ( .A1(G85), .A2(n649), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U712 ( .A(KEYINPUT66), .B(n635), .Z(n639) );
  NAND2_X1 U713 ( .A1(G60), .A2(n660), .ZN(n637) );
  NAND2_X1 U714 ( .A1(G47), .A2(n656), .ZN(n636) );
  AND2_X1 U715 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(G290) );
  NAND2_X1 U717 ( .A1(G48), .A2(n656), .ZN(n640) );
  XNOR2_X1 U718 ( .A(n640), .B(KEYINPUT80), .ZN(n647) );
  NAND2_X1 U719 ( .A1(n660), .A2(G61), .ZN(n642) );
  NAND2_X1 U720 ( .A1(G86), .A2(n649), .ZN(n641) );
  NAND2_X1 U721 ( .A1(n642), .A2(n641), .ZN(n645) );
  NAND2_X1 U722 ( .A1(n648), .A2(G73), .ZN(n643) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n643), .Z(n644) );
  NOR2_X1 U724 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n647), .A2(n646), .ZN(G305) );
  NAND2_X1 U726 ( .A1(n648), .A2(G75), .ZN(n651) );
  NAND2_X1 U727 ( .A1(G88), .A2(n649), .ZN(n650) );
  NAND2_X1 U728 ( .A1(n651), .A2(n650), .ZN(n655) );
  NAND2_X1 U729 ( .A1(G62), .A2(n660), .ZN(n653) );
  NAND2_X1 U730 ( .A1(G50), .A2(n656), .ZN(n652) );
  NAND2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U732 ( .A1(n655), .A2(n654), .ZN(G166) );
  NAND2_X1 U733 ( .A1(G49), .A2(n656), .ZN(n658) );
  NAND2_X1 U734 ( .A1(G74), .A2(G651), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U736 ( .A1(n660), .A2(n659), .ZN(n664) );
  NAND2_X1 U737 ( .A1(G87), .A2(n661), .ZN(n662) );
  XOR2_X1 U738 ( .A(KEYINPUT79), .B(n662), .Z(n663) );
  NAND2_X1 U739 ( .A1(n664), .A2(n663), .ZN(G288) );
  XNOR2_X1 U740 ( .A(G290), .B(G305), .ZN(n670) );
  XOR2_X1 U741 ( .A(KEYINPUT81), .B(KEYINPUT19), .Z(n666) );
  XNOR2_X1 U742 ( .A(G166), .B(KEYINPUT82), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U744 ( .A(n674), .B(n667), .ZN(n668) );
  XNOR2_X1 U745 ( .A(n668), .B(G288), .ZN(n669) );
  XNOR2_X1 U746 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U747 ( .A(G299), .B(n671), .ZN(n893) );
  XNOR2_X1 U748 ( .A(n672), .B(n893), .ZN(n673) );
  NAND2_X1 U749 ( .A1(n673), .A2(G868), .ZN(n676) );
  OR2_X1 U750 ( .A1(G868), .A2(n674), .ZN(n675) );
  NAND2_X1 U751 ( .A1(n676), .A2(n675), .ZN(G295) );
  NAND2_X1 U752 ( .A1(G2078), .A2(G2084), .ZN(n677) );
  XOR2_X1 U753 ( .A(KEYINPUT20), .B(n677), .Z(n678) );
  NAND2_X1 U754 ( .A1(G2090), .A2(n678), .ZN(n679) );
  XNOR2_X1 U755 ( .A(KEYINPUT21), .B(n679), .ZN(n680) );
  NAND2_X1 U756 ( .A1(n680), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U757 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U758 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NAND2_X1 U759 ( .A1(G661), .A2(G483), .ZN(n689) );
  NOR2_X1 U760 ( .A1(G219), .A2(G220), .ZN(n681) );
  XOR2_X1 U761 ( .A(KEYINPUT22), .B(n681), .Z(n682) );
  NOR2_X1 U762 ( .A1(G218), .A2(n682), .ZN(n683) );
  XOR2_X1 U763 ( .A(KEYINPUT83), .B(n683), .Z(n684) );
  NAND2_X1 U764 ( .A1(G96), .A2(n684), .ZN(n846) );
  NAND2_X1 U765 ( .A1(n846), .A2(G2106), .ZN(n688) );
  NAND2_X1 U766 ( .A1(G69), .A2(G120), .ZN(n685) );
  NOR2_X1 U767 ( .A1(G237), .A2(n685), .ZN(n686) );
  NAND2_X1 U768 ( .A1(G108), .A2(n686), .ZN(n847) );
  NAND2_X1 U769 ( .A1(n847), .A2(G567), .ZN(n687) );
  NAND2_X1 U770 ( .A1(n688), .A2(n687), .ZN(n924) );
  NOR2_X1 U771 ( .A1(n689), .A2(n924), .ZN(n690) );
  XNOR2_X1 U772 ( .A(n690), .B(KEYINPUT84), .ZN(n845) );
  NAND2_X1 U773 ( .A1(G36), .A2(n845), .ZN(G176) );
  INV_X1 U774 ( .A(G166), .ZN(G303) );
  NOR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n796) );
  INV_X1 U776 ( .A(G40), .ZN(n691) );
  OR2_X1 U777 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U778 ( .A1(n694), .A2(n693), .ZN(n794) );
  AND2_X1 U779 ( .A1(n796), .A2(n794), .ZN(n729) );
  NAND2_X1 U780 ( .A1(G8), .A2(n744), .ZN(n773) );
  NOR2_X1 U781 ( .A1(G1981), .A2(G305), .ZN(n695) );
  XOR2_X1 U782 ( .A(n695), .B(KEYINPUT24), .Z(n696) );
  NOR2_X1 U783 ( .A1(n773), .A2(n696), .ZN(n783) );
  AND2_X1 U784 ( .A1(n951), .A2(n697), .ZN(n702) );
  NAND2_X1 U785 ( .A1(G1996), .A2(n729), .ZN(n698) );
  XNOR2_X1 U786 ( .A(n698), .B(KEYINPUT26), .ZN(n700) );
  NAND2_X1 U787 ( .A1(G1341), .A2(n744), .ZN(n699) );
  NAND2_X1 U788 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U789 ( .A(KEYINPUT95), .B(n701), .ZN(n713) );
  AND2_X1 U790 ( .A1(n702), .A2(n713), .ZN(n703) );
  XOR2_X1 U791 ( .A(n703), .B(KEYINPUT96), .Z(n712) );
  NAND2_X1 U792 ( .A1(G2067), .A2(n729), .ZN(n704) );
  XNOR2_X1 U793 ( .A(KEYINPUT98), .B(n704), .ZN(n705) );
  NAND2_X1 U794 ( .A1(n744), .A2(G1348), .ZN(n707) );
  NAND2_X1 U795 ( .A1(n705), .A2(n707), .ZN(n706) );
  NOR2_X1 U796 ( .A1(KEYINPUT97), .A2(n706), .ZN(n710) );
  NAND2_X1 U797 ( .A1(KEYINPUT98), .A2(KEYINPUT97), .ZN(n708) );
  NOR2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U799 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U800 ( .A1(n712), .A2(n711), .ZN(n721) );
  NAND2_X1 U801 ( .A1(n713), .A2(n951), .ZN(n714) );
  NAND2_X1 U802 ( .A1(n714), .A2(n952), .ZN(n719) );
  NAND2_X1 U803 ( .A1(n729), .A2(G2072), .ZN(n715) );
  XNOR2_X1 U804 ( .A(n715), .B(KEYINPUT27), .ZN(n717) );
  INV_X1 U805 ( .A(G1956), .ZN(n975) );
  NOR2_X1 U806 ( .A1(n975), .A2(n729), .ZN(n716) );
  NOR2_X1 U807 ( .A1(n717), .A2(n716), .ZN(n723) );
  NOR2_X1 U808 ( .A1(n955), .A2(n723), .ZN(n718) );
  XOR2_X1 U809 ( .A(n718), .B(KEYINPUT28), .Z(n722) );
  AND2_X1 U810 ( .A1(n719), .A2(n722), .ZN(n720) );
  NAND2_X1 U811 ( .A1(n721), .A2(n720), .ZN(n727) );
  INV_X1 U812 ( .A(n722), .ZN(n725) );
  NAND2_X1 U813 ( .A1(n955), .A2(n723), .ZN(n724) );
  OR2_X1 U814 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U815 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U816 ( .A(n728), .B(KEYINPUT29), .ZN(n733) );
  XNOR2_X1 U817 ( .A(G2078), .B(KEYINPUT25), .ZN(n936) );
  NOR2_X1 U818 ( .A1(n744), .A2(n936), .ZN(n731) );
  INV_X1 U819 ( .A(G1961), .ZN(n974) );
  NOR2_X1 U820 ( .A1(n729), .A2(n974), .ZN(n730) );
  NOR2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n737) );
  NAND2_X1 U822 ( .A1(G171), .A2(n737), .ZN(n732) );
  NAND2_X1 U823 ( .A1(n733), .A2(n732), .ZN(n743) );
  NOR2_X1 U824 ( .A1(G1966), .A2(n773), .ZN(n755) );
  NOR2_X1 U825 ( .A1(G2084), .A2(n744), .ZN(n752) );
  NOR2_X1 U826 ( .A1(n755), .A2(n752), .ZN(n734) );
  NAND2_X1 U827 ( .A1(G8), .A2(n734), .ZN(n735) );
  XNOR2_X1 U828 ( .A(KEYINPUT30), .B(n735), .ZN(n736) );
  NOR2_X1 U829 ( .A1(G168), .A2(n736), .ZN(n739) );
  NOR2_X1 U830 ( .A1(G171), .A2(n737), .ZN(n738) );
  NOR2_X1 U831 ( .A1(n739), .A2(n738), .ZN(n741) );
  NAND2_X1 U832 ( .A1(n743), .A2(n742), .ZN(n753) );
  NAND2_X1 U833 ( .A1(n753), .A2(G286), .ZN(n749) );
  NOR2_X1 U834 ( .A1(G1971), .A2(n773), .ZN(n746) );
  NOR2_X1 U835 ( .A1(G2090), .A2(n744), .ZN(n745) );
  NOR2_X1 U836 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U837 ( .A1(n747), .A2(G303), .ZN(n748) );
  NAND2_X1 U838 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U839 ( .A1(G8), .A2(n750), .ZN(n751) );
  XNOR2_X1 U840 ( .A(KEYINPUT32), .B(n751), .ZN(n759) );
  NAND2_X1 U841 ( .A1(G8), .A2(n752), .ZN(n757) );
  INV_X1 U842 ( .A(n753), .ZN(n754) );
  NOR2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U844 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U845 ( .A1(n759), .A2(n758), .ZN(n765) );
  NOR2_X1 U846 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U847 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n765), .A2(n761), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n762), .A2(n773), .ZN(n781) );
  NOR2_X1 U850 ( .A1(G1976), .A2(G288), .ZN(n768) );
  NOR2_X1 U851 ( .A1(G1971), .A2(G303), .ZN(n763) );
  NOR2_X1 U852 ( .A1(n768), .A2(n763), .ZN(n959) );
  XNOR2_X1 U853 ( .A(KEYINPUT100), .B(n959), .ZN(n764) );
  NAND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n766) );
  NAND2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n958) );
  NAND2_X1 U856 ( .A1(n766), .A2(n958), .ZN(n775) );
  XOR2_X1 U857 ( .A(G1981), .B(KEYINPUT102), .Z(n767) );
  XNOR2_X1 U858 ( .A(G305), .B(n767), .ZN(n948) );
  INV_X1 U859 ( .A(n948), .ZN(n772) );
  NAND2_X1 U860 ( .A1(KEYINPUT33), .A2(n768), .ZN(n769) );
  XOR2_X1 U861 ( .A(KEYINPUT101), .B(n769), .Z(n770) );
  NOR2_X1 U862 ( .A1(n773), .A2(n770), .ZN(n771) );
  OR2_X1 U863 ( .A1(n772), .A2(n771), .ZN(n776) );
  OR2_X1 U864 ( .A1(n773), .A2(n776), .ZN(n774) );
  NOR2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n779) );
  INV_X1 U866 ( .A(n776), .ZN(n777) );
  AND2_X1 U867 ( .A1(n777), .A2(KEYINPUT33), .ZN(n778) );
  NOR2_X1 U868 ( .A1(n779), .A2(n778), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U870 ( .A1(n783), .A2(n526), .ZN(n823) );
  XNOR2_X1 U871 ( .A(KEYINPUT37), .B(G2067), .ZN(n834) );
  NAND2_X1 U872 ( .A1(n873), .A2(G128), .ZN(n784) );
  XNOR2_X1 U873 ( .A(n784), .B(KEYINPUT88), .ZN(n786) );
  NAND2_X1 U874 ( .A1(G116), .A2(n874), .ZN(n785) );
  NAND2_X1 U875 ( .A1(n786), .A2(n785), .ZN(n787) );
  XNOR2_X1 U876 ( .A(n787), .B(KEYINPUT35), .ZN(n792) );
  NAND2_X1 U877 ( .A1(G140), .A2(n869), .ZN(n789) );
  NAND2_X1 U878 ( .A1(G104), .A2(n870), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U880 ( .A(KEYINPUT34), .B(n790), .Z(n791) );
  NAND2_X1 U881 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U882 ( .A(n793), .B(KEYINPUT36), .Z(n888) );
  OR2_X1 U883 ( .A1(n834), .A2(n888), .ZN(n1015) );
  INV_X1 U884 ( .A(n794), .ZN(n795) );
  NOR2_X1 U885 ( .A1(n796), .A2(n795), .ZN(n797) );
  XOR2_X1 U886 ( .A(KEYINPUT87), .B(n797), .Z(n836) );
  INV_X1 U887 ( .A(n836), .ZN(n818) );
  NOR2_X1 U888 ( .A1(n1015), .A2(n818), .ZN(n798) );
  XNOR2_X1 U889 ( .A(n798), .B(KEYINPUT89), .ZN(n831) );
  NAND2_X1 U890 ( .A1(G129), .A2(n873), .ZN(n800) );
  NAND2_X1 U891 ( .A1(G117), .A2(n874), .ZN(n799) );
  NAND2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n801) );
  XNOR2_X1 U893 ( .A(KEYINPUT92), .B(n801), .ZN(n804) );
  NAND2_X1 U894 ( .A1(n870), .A2(G105), .ZN(n802) );
  XOR2_X1 U895 ( .A(KEYINPUT38), .B(n802), .Z(n803) );
  NOR2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n806) );
  NAND2_X1 U897 ( .A1(n869), .A2(G141), .ZN(n805) );
  NAND2_X1 U898 ( .A1(n806), .A2(n805), .ZN(n864) );
  NAND2_X1 U899 ( .A1(n864), .A2(G1996), .ZN(n816) );
  NAND2_X1 U900 ( .A1(G107), .A2(n874), .ZN(n807) );
  XOR2_X1 U901 ( .A(KEYINPUT90), .B(n807), .Z(n812) );
  NAND2_X1 U902 ( .A1(G131), .A2(n869), .ZN(n809) );
  NAND2_X1 U903 ( .A1(G95), .A2(n870), .ZN(n808) );
  NAND2_X1 U904 ( .A1(n809), .A2(n808), .ZN(n810) );
  XOR2_X1 U905 ( .A(KEYINPUT91), .B(n810), .Z(n811) );
  NOR2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U907 ( .A1(n873), .A2(G119), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n814), .A2(n813), .ZN(n865) );
  NAND2_X1 U909 ( .A1(G1991), .A2(n865), .ZN(n815) );
  NAND2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U911 ( .A(n817), .B(KEYINPUT93), .ZN(n1024) );
  XNOR2_X1 U912 ( .A(KEYINPUT94), .B(n818), .ZN(n819) );
  NOR2_X1 U913 ( .A1(n1024), .A2(n819), .ZN(n827) );
  INV_X1 U914 ( .A(n827), .ZN(n820) );
  NAND2_X1 U915 ( .A1(n831), .A2(n820), .ZN(n822) );
  XNOR2_X1 U916 ( .A(G1986), .B(KEYINPUT86), .ZN(n821) );
  XNOR2_X1 U917 ( .A(n821), .B(G290), .ZN(n954) );
  NOR2_X1 U918 ( .A1(n864), .A2(G1996), .ZN(n824) );
  XNOR2_X1 U919 ( .A(n824), .B(KEYINPUT104), .ZN(n1007) );
  NOR2_X1 U920 ( .A1(G1991), .A2(n865), .ZN(n1014) );
  NOR2_X1 U921 ( .A1(G1986), .A2(G290), .ZN(n825) );
  NOR2_X1 U922 ( .A1(n1014), .A2(n825), .ZN(n826) );
  NOR2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  XOR2_X1 U924 ( .A(KEYINPUT105), .B(n828), .Z(n829) );
  NOR2_X1 U925 ( .A1(n1007), .A2(n829), .ZN(n830) );
  XNOR2_X1 U926 ( .A(n830), .B(KEYINPUT39), .ZN(n832) );
  NAND2_X1 U927 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U928 ( .A(n833), .B(KEYINPUT106), .ZN(n835) );
  NAND2_X1 U929 ( .A1(n834), .A2(n888), .ZN(n1009) );
  NAND2_X1 U930 ( .A1(n835), .A2(n1009), .ZN(n837) );
  NAND2_X1 U931 ( .A1(n837), .A2(n836), .ZN(n838) );
  NAND2_X1 U932 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U933 ( .A(KEYINPUT40), .B(n840), .ZN(G329) );
  NAND2_X1 U934 ( .A1(n841), .A2(G2106), .ZN(n842) );
  XNOR2_X1 U935 ( .A(n842), .B(KEYINPUT108), .ZN(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n843) );
  NAND2_X1 U937 ( .A1(G661), .A2(n843), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n844) );
  NAND2_X1 U939 ( .A1(n845), .A2(n844), .ZN(G188) );
  INV_X1 U941 ( .A(G120), .ZN(G236) );
  INV_X1 U942 ( .A(G96), .ZN(G221) );
  INV_X1 U943 ( .A(G69), .ZN(G235) );
  NOR2_X1 U944 ( .A1(n847), .A2(n846), .ZN(G325) );
  INV_X1 U945 ( .A(G325), .ZN(G261) );
  NAND2_X1 U946 ( .A1(n873), .A2(G124), .ZN(n848) );
  XNOR2_X1 U947 ( .A(n848), .B(KEYINPUT44), .ZN(n850) );
  NAND2_X1 U948 ( .A1(G112), .A2(n874), .ZN(n849) );
  NAND2_X1 U949 ( .A1(n850), .A2(n849), .ZN(n854) );
  NAND2_X1 U950 ( .A1(G136), .A2(n869), .ZN(n852) );
  NAND2_X1 U951 ( .A1(G100), .A2(n870), .ZN(n851) );
  NAND2_X1 U952 ( .A1(n852), .A2(n851), .ZN(n853) );
  NOR2_X1 U953 ( .A1(n854), .A2(n853), .ZN(G162) );
  NAND2_X1 U954 ( .A1(n870), .A2(G106), .ZN(n855) );
  XOR2_X1 U955 ( .A(KEYINPUT113), .B(n855), .Z(n857) );
  NAND2_X1 U956 ( .A1(n869), .A2(G142), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n858), .B(KEYINPUT45), .ZN(n860) );
  NAND2_X1 U959 ( .A1(G118), .A2(n874), .ZN(n859) );
  NAND2_X1 U960 ( .A1(n860), .A2(n859), .ZN(n863) );
  NAND2_X1 U961 ( .A1(n873), .A2(G130), .ZN(n861) );
  XOR2_X1 U962 ( .A(KEYINPUT112), .B(n861), .Z(n862) );
  NOR2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n868) );
  XNOR2_X1 U964 ( .A(G162), .B(n864), .ZN(n866) );
  XNOR2_X1 U965 ( .A(n866), .B(n865), .ZN(n867) );
  XOR2_X1 U966 ( .A(n868), .B(n867), .Z(n881) );
  NAND2_X1 U967 ( .A1(G139), .A2(n869), .ZN(n872) );
  NAND2_X1 U968 ( .A1(G103), .A2(n870), .ZN(n871) );
  NAND2_X1 U969 ( .A1(n872), .A2(n871), .ZN(n879) );
  NAND2_X1 U970 ( .A1(G127), .A2(n873), .ZN(n876) );
  NAND2_X1 U971 ( .A1(G115), .A2(n874), .ZN(n875) );
  NAND2_X1 U972 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U973 ( .A(KEYINPUT47), .B(n877), .Z(n878) );
  NOR2_X1 U974 ( .A1(n879), .A2(n878), .ZN(n1017) );
  XNOR2_X1 U975 ( .A(G160), .B(n1017), .ZN(n880) );
  XNOR2_X1 U976 ( .A(n881), .B(n880), .ZN(n890) );
  XNOR2_X1 U977 ( .A(KEYINPUT116), .B(KEYINPUT48), .ZN(n883) );
  XNOR2_X1 U978 ( .A(n1011), .B(KEYINPUT115), .ZN(n882) );
  XNOR2_X1 U979 ( .A(n883), .B(n882), .ZN(n884) );
  XOR2_X1 U980 ( .A(n884), .B(KEYINPUT46), .Z(n886) );
  XNOR2_X1 U981 ( .A(G164), .B(KEYINPUT114), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U983 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U984 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U985 ( .A1(G37), .A2(n891), .ZN(G395) );
  XNOR2_X1 U986 ( .A(G171), .B(n952), .ZN(n892) );
  XNOR2_X1 U987 ( .A(n892), .B(G286), .ZN(n895) );
  XNOR2_X1 U988 ( .A(n951), .B(n893), .ZN(n894) );
  XNOR2_X1 U989 ( .A(n895), .B(n894), .ZN(n896) );
  NOR2_X1 U990 ( .A1(G37), .A2(n896), .ZN(G397) );
  XOR2_X1 U991 ( .A(KEYINPUT42), .B(G2084), .Z(n898) );
  XNOR2_X1 U992 ( .A(G2078), .B(G2072), .ZN(n897) );
  XNOR2_X1 U993 ( .A(n898), .B(n897), .ZN(n899) );
  XOR2_X1 U994 ( .A(n899), .B(G2096), .Z(n901) );
  XNOR2_X1 U995 ( .A(G2067), .B(G2090), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n901), .B(n900), .ZN(n905) );
  XOR2_X1 U997 ( .A(KEYINPUT43), .B(G2678), .Z(n903) );
  XNOR2_X1 U998 ( .A(KEYINPUT109), .B(G2100), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1000 ( .A(n905), .B(n904), .Z(G227) );
  XOR2_X1 U1001 ( .A(KEYINPUT41), .B(G1961), .Z(n907) );
  XNOR2_X1 U1002 ( .A(G1981), .B(G1966), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1004 ( .A(n908), .B(G2474), .Z(n910) );
  XNOR2_X1 U1005 ( .A(G1996), .B(G1991), .ZN(n909) );
  XNOR2_X1 U1006 ( .A(n910), .B(n909), .ZN(n914) );
  XOR2_X1 U1007 ( .A(G1971), .B(G1956), .Z(n912) );
  XNOR2_X1 U1008 ( .A(G1986), .B(G1976), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n912), .B(n911), .ZN(n913) );
  XOR2_X1 U1010 ( .A(n914), .B(n913), .Z(n916) );
  XNOR2_X1 U1011 ( .A(KEYINPUT111), .B(KEYINPUT110), .ZN(n915) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(G229) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1014 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1015 ( .A1(G397), .A2(n918), .ZN(n921) );
  NOR2_X1 U1016 ( .A1(n924), .A2(G401), .ZN(n919) );
  XOR2_X1 U1017 ( .A(KEYINPUT117), .B(n919), .Z(n920) );
  NAND2_X1 U1018 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1019 ( .A1(G395), .A2(n922), .ZN(n923) );
  XNOR2_X1 U1020 ( .A(KEYINPUT118), .B(n923), .ZN(G308) );
  INV_X1 U1021 ( .A(G308), .ZN(G225) );
  INV_X1 U1022 ( .A(n924), .ZN(G319) );
  INV_X1 U1023 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1024 ( .A(G2090), .B(KEYINPUT119), .ZN(n925) );
  XNOR2_X1 U1025 ( .A(n925), .B(G35), .ZN(n928) );
  XOR2_X1 U1026 ( .A(G2084), .B(G34), .Z(n926) );
  XNOR2_X1 U1027 ( .A(KEYINPUT54), .B(n926), .ZN(n927) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n942) );
  XNOR2_X1 U1029 ( .A(G2067), .B(G26), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(G33), .B(G2072), .ZN(n929) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n935) );
  XOR2_X1 U1032 ( .A(G1991), .B(G25), .Z(n931) );
  NAND2_X1 U1033 ( .A1(n931), .A2(G28), .ZN(n933) );
  XNOR2_X1 U1034 ( .A(G32), .B(G1996), .ZN(n932) );
  NOR2_X1 U1035 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1036 ( .A1(n935), .A2(n934), .ZN(n938) );
  XOR2_X1 U1037 ( .A(G27), .B(n936), .Z(n937) );
  NOR2_X1 U1038 ( .A1(n938), .A2(n937), .ZN(n939) );
  XNOR2_X1 U1039 ( .A(KEYINPUT120), .B(n939), .ZN(n940) );
  XNOR2_X1 U1040 ( .A(KEYINPUT53), .B(n940), .ZN(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1042 ( .A(KEYINPUT55), .B(n943), .ZN(n945) );
  INV_X1 U1043 ( .A(G29), .ZN(n944) );
  NAND2_X1 U1044 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1045 ( .A1(n946), .A2(G11), .ZN(n947) );
  XNOR2_X1 U1046 ( .A(KEYINPUT121), .B(n947), .ZN(n1004) );
  XNOR2_X1 U1047 ( .A(G16), .B(KEYINPUT56), .ZN(n973) );
  XNOR2_X1 U1048 ( .A(G1966), .B(G168), .ZN(n949) );
  NAND2_X1 U1049 ( .A1(n949), .A2(n948), .ZN(n950) );
  XNOR2_X1 U1050 ( .A(n950), .B(KEYINPUT57), .ZN(n971) );
  XOR2_X1 U1051 ( .A(n951), .B(G1341), .Z(n969) );
  XNOR2_X1 U1052 ( .A(G1348), .B(n952), .ZN(n953) );
  NOR2_X1 U1053 ( .A1(n954), .A2(n953), .ZN(n964) );
  XNOR2_X1 U1054 ( .A(n955), .B(G1956), .ZN(n957) );
  NAND2_X1 U1055 ( .A1(G1971), .A2(G303), .ZN(n956) );
  NAND2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n961) );
  NAND2_X1 U1057 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1059 ( .A(n962), .B(KEYINPUT122), .ZN(n963) );
  NAND2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n966) );
  XNOR2_X1 U1061 ( .A(G1961), .B(G301), .ZN(n965) );
  NOR2_X1 U1062 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1063 ( .A(KEYINPUT123), .B(n967), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n1001) );
  INV_X1 U1067 ( .A(G16), .ZN(n999) );
  XNOR2_X1 U1068 ( .A(n974), .B(G5), .ZN(n995) );
  XOR2_X1 U1069 ( .A(G1966), .B(G21), .Z(n985) );
  XNOR2_X1 U1070 ( .A(G20), .B(n975), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(G1981), .B(G6), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(G19), .B(G1341), .ZN(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n982) );
  XOR2_X1 U1075 ( .A(KEYINPUT59), .B(G1348), .Z(n980) );
  XNOR2_X1 U1076 ( .A(G4), .B(n980), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1078 ( .A(n983), .B(KEYINPUT60), .ZN(n984) );
  NAND2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n986) );
  XNOR2_X1 U1080 ( .A(KEYINPUT124), .B(n986), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(G1976), .B(G23), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(G1971), .B(G22), .ZN(n987) );
  NOR2_X1 U1083 ( .A1(n988), .A2(n987), .ZN(n990) );
  XOR2_X1 U1084 ( .A(G1986), .B(G24), .Z(n989) );
  NAND2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1086 ( .A(KEYINPUT58), .B(n991), .ZN(n992) );
  NOR2_X1 U1087 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1088 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1089 ( .A(n996), .B(KEYINPUT61), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(KEYINPUT125), .B(n997), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1093 ( .A(KEYINPUT126), .B(n1002), .Z(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XNOR2_X1 U1095 ( .A(n1005), .B(KEYINPUT127), .ZN(n1032) );
  XOR2_X1 U1096 ( .A(G2090), .B(G162), .Z(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1098 ( .A(KEYINPUT51), .B(n1008), .Z(n1010) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1026) );
  XNOR2_X1 U1100 ( .A(G160), .B(G2084), .ZN(n1012) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1022) );
  XOR2_X1 U1104 ( .A(G2072), .B(n1017), .Z(n1019) );
  XOR2_X1 U1105 ( .A(G164), .B(G2078), .Z(n1018) );
  NOR2_X1 U1106 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1107 ( .A(KEYINPUT50), .B(n1020), .Z(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(KEYINPUT52), .B(n1027), .ZN(n1029) );
  INV_X1 U1112 ( .A(KEYINPUT55), .ZN(n1028) );
  NAND2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(n1030), .A2(G29), .ZN(n1031) );
  NAND2_X1 U1115 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1033), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

