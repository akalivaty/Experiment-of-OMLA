

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578;

  NOR2_X2 U318 ( .A1(n524), .A2(n441), .ZN(n442) );
  XOR2_X1 U319 ( .A(KEYINPUT119), .B(n442), .Z(n553) );
  XOR2_X1 U320 ( .A(n350), .B(n349), .Z(n549) );
  AND2_X1 U321 ( .A1(G232GAT), .A2(G233GAT), .ZN(n286) );
  XNOR2_X1 U322 ( .A(n394), .B(KEYINPUT47), .ZN(n395) );
  XNOR2_X1 U323 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U324 ( .A(n349), .B(n332), .ZN(n333) );
  XNOR2_X1 U325 ( .A(n345), .B(n286), .ZN(n346) );
  XNOR2_X1 U326 ( .A(n334), .B(n333), .ZN(n389) );
  XNOR2_X1 U327 ( .A(n347), .B(n346), .ZN(n348) );
  INV_X1 U328 ( .A(n540), .ZN(n526) );
  XNOR2_X1 U329 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n444) );
  XNOR2_X1 U330 ( .A(n445), .B(n444), .ZN(G1351GAT) );
  XOR2_X1 U331 ( .A(G176GAT), .B(KEYINPUT83), .Z(n288) );
  XNOR2_X1 U332 ( .A(G169GAT), .B(KEYINPUT84), .ZN(n287) );
  XNOR2_X1 U333 ( .A(n288), .B(n287), .ZN(n305) );
  XOR2_X1 U334 ( .A(G134GAT), .B(G99GAT), .Z(n290) );
  XNOR2_X1 U335 ( .A(G43GAT), .B(G190GAT), .ZN(n289) );
  XNOR2_X1 U336 ( .A(n290), .B(n289), .ZN(n294) );
  XOR2_X1 U337 ( .A(KEYINPUT20), .B(G120GAT), .Z(n292) );
  XNOR2_X1 U338 ( .A(G113GAT), .B(G15GAT), .ZN(n291) );
  XNOR2_X1 U339 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U340 ( .A(n294), .B(n293), .Z(n303) );
  XOR2_X1 U341 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n296) );
  XNOR2_X1 U342 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n295) );
  XNOR2_X1 U343 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U344 ( .A(KEYINPUT19), .B(n297), .Z(n306) );
  XNOR2_X1 U345 ( .A(G127GAT), .B(KEYINPUT81), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n298), .B(KEYINPUT0), .ZN(n408) );
  XOR2_X1 U347 ( .A(n408), .B(G71GAT), .Z(n300) );
  NAND2_X1 U348 ( .A1(G227GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U349 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n306), .B(n301), .ZN(n302) );
  XNOR2_X1 U351 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U352 ( .A(n305), .B(n304), .Z(n524) );
  XOR2_X1 U353 ( .A(G190GAT), .B(G218GAT), .Z(n340) );
  XOR2_X1 U354 ( .A(G176GAT), .B(G64GAT), .Z(n331) );
  XOR2_X1 U355 ( .A(n331), .B(G92GAT), .Z(n308) );
  XNOR2_X1 U356 ( .A(G36GAT), .B(n306), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U358 ( .A(n340), .B(n309), .Z(n313) );
  XOR2_X1 U359 ( .A(G169GAT), .B(G8GAT), .Z(n385) );
  XOR2_X1 U360 ( .A(G204GAT), .B(G211GAT), .Z(n311) );
  XNOR2_X1 U361 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n426) );
  XNOR2_X1 U363 ( .A(n385), .B(n426), .ZN(n312) );
  XNOR2_X1 U364 ( .A(n313), .B(n312), .ZN(n318) );
  XOR2_X1 U365 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n315) );
  NAND2_X1 U366 ( .A1(G226GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U368 ( .A(KEYINPUT92), .B(n316), .Z(n317) );
  XNOR2_X1 U369 ( .A(n318), .B(n317), .ZN(n472) );
  XOR2_X1 U370 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n320) );
  NAND2_X1 U371 ( .A1(G230GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U372 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U373 ( .A(n321), .B(KEYINPUT31), .Z(n326) );
  XOR2_X1 U374 ( .A(KEYINPUT71), .B(KEYINPUT13), .Z(n323) );
  XNOR2_X1 U375 ( .A(G71GAT), .B(G78GAT), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n360) );
  XNOR2_X1 U377 ( .A(G120GAT), .B(G148GAT), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n324), .B(G57GAT), .ZN(n407) );
  XNOR2_X1 U379 ( .A(n360), .B(n407), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n326), .B(n325), .ZN(n327) );
  XOR2_X1 U381 ( .A(n327), .B(KEYINPUT32), .Z(n334) );
  XOR2_X1 U382 ( .A(KEYINPUT73), .B(G92GAT), .Z(n329) );
  XNOR2_X1 U383 ( .A(G99GAT), .B(G106GAT), .ZN(n328) );
  XNOR2_X1 U384 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U385 ( .A(G85GAT), .B(n330), .ZN(n349) );
  XNOR2_X1 U386 ( .A(G204GAT), .B(n331), .ZN(n332) );
  XOR2_X1 U387 ( .A(G43GAT), .B(G29GAT), .Z(n336) );
  XNOR2_X1 U388 ( .A(G50GAT), .B(KEYINPUT8), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U390 ( .A(n337), .B(KEYINPUT7), .Z(n339) );
  XNOR2_X1 U391 ( .A(G36GAT), .B(KEYINPUT66), .ZN(n338) );
  XNOR2_X1 U392 ( .A(n339), .B(n338), .ZN(n380) );
  XOR2_X1 U393 ( .A(KEYINPUT10), .B(KEYINPUT74), .Z(n342) );
  XOR2_X1 U394 ( .A(G134GAT), .B(G162GAT), .Z(n411) );
  XNOR2_X1 U395 ( .A(n411), .B(n340), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n347) );
  XOR2_X1 U397 ( .A(KEYINPUT75), .B(KEYINPUT76), .Z(n344) );
  XNOR2_X1 U398 ( .A(KEYINPUT9), .B(KEYINPUT11), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n345) );
  XNOR2_X1 U400 ( .A(n380), .B(n348), .ZN(n350) );
  XNOR2_X1 U401 ( .A(KEYINPUT77), .B(n549), .ZN(n443) );
  XOR2_X1 U402 ( .A(KEYINPUT36), .B(n443), .Z(n575) );
  XOR2_X1 U403 ( .A(KEYINPUT12), .B(KEYINPUT15), .Z(n352) );
  XNOR2_X1 U404 ( .A(G8GAT), .B(G64GAT), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n352), .B(n351), .ZN(n368) );
  XOR2_X1 U406 ( .A(G57GAT), .B(G127GAT), .Z(n354) );
  XNOR2_X1 U407 ( .A(G1GAT), .B(G183GAT), .ZN(n353) );
  XNOR2_X1 U408 ( .A(n354), .B(n353), .ZN(n356) );
  XOR2_X1 U409 ( .A(G155GAT), .B(G211GAT), .Z(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n364) );
  XNOR2_X1 U411 ( .A(KEYINPUT78), .B(KEYINPUT80), .ZN(n357) );
  XNOR2_X1 U412 ( .A(n357), .B(KEYINPUT79), .ZN(n358) );
  XOR2_X1 U413 ( .A(n358), .B(KEYINPUT14), .Z(n362) );
  XNOR2_X1 U414 ( .A(G22GAT), .B(G15GAT), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n359), .B(KEYINPUT67), .ZN(n383) );
  XNOR2_X1 U416 ( .A(n383), .B(n360), .ZN(n361) );
  XNOR2_X1 U417 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U418 ( .A(n364), .B(n363), .ZN(n366) );
  NAND2_X1 U419 ( .A1(G231GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U421 ( .A(n368), .B(n367), .ZN(n544) );
  NOR2_X1 U422 ( .A1(n575), .A2(n544), .ZN(n370) );
  INV_X1 U423 ( .A(KEYINPUT45), .ZN(n369) );
  XNOR2_X1 U424 ( .A(n370), .B(n369), .ZN(n371) );
  NOR2_X1 U425 ( .A1(n389), .A2(n371), .ZN(n373) );
  INV_X1 U426 ( .A(KEYINPUT112), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n388) );
  XOR2_X1 U428 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n375) );
  NAND2_X1 U429 ( .A1(G229GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U430 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U431 ( .A(n376), .B(KEYINPUT69), .Z(n382) );
  XOR2_X1 U432 ( .A(KEYINPUT68), .B(KEYINPUT29), .Z(n378) );
  XNOR2_X1 U433 ( .A(G141GAT), .B(G197GAT), .ZN(n377) );
  XNOR2_X1 U434 ( .A(n378), .B(n377), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n384) );
  XOR2_X1 U437 ( .A(n384), .B(n383), .Z(n387) );
  XOR2_X1 U438 ( .A(G113GAT), .B(G1GAT), .Z(n412) );
  XNOR2_X1 U439 ( .A(n412), .B(n385), .ZN(n386) );
  XNOR2_X1 U440 ( .A(n387), .B(n386), .ZN(n563) );
  XNOR2_X1 U441 ( .A(KEYINPUT70), .B(n563), .ZN(n551) );
  NOR2_X1 U442 ( .A1(n388), .A2(n551), .ZN(n398) );
  INV_X1 U443 ( .A(n544), .ZN(n570) );
  INV_X1 U444 ( .A(n389), .ZN(n450) );
  XOR2_X1 U445 ( .A(KEYINPUT41), .B(n450), .Z(n540) );
  NAND2_X1 U446 ( .A1(n526), .A2(n563), .ZN(n391) );
  XOR2_X1 U447 ( .A(KEYINPUT109), .B(KEYINPUT46), .Z(n390) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n392) );
  NAND2_X1 U449 ( .A1(n392), .A2(n549), .ZN(n393) );
  NOR2_X1 U450 ( .A1(n570), .A2(n393), .ZN(n396) );
  XNOR2_X1 U451 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n394) );
  NOR2_X1 U452 ( .A1(n398), .A2(n397), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n399), .B(KEYINPUT48), .ZN(n521) );
  NOR2_X1 U454 ( .A1(n472), .A2(n521), .ZN(n400) );
  XNOR2_X1 U455 ( .A(n400), .B(KEYINPUT54), .ZN(n559) );
  XOR2_X1 U456 ( .A(KEYINPUT3), .B(KEYINPUT86), .Z(n402) );
  XNOR2_X1 U457 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n401) );
  XNOR2_X1 U458 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U459 ( .A(G141GAT), .B(n403), .Z(n433) );
  XOR2_X1 U460 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n405) );
  NAND2_X1 U461 ( .A1(G225GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U462 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U463 ( .A(n406), .B(KEYINPUT1), .Z(n410) );
  XNOR2_X1 U464 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U465 ( .A(n410), .B(n409), .ZN(n416) );
  XOR2_X1 U466 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n414) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U468 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U469 ( .A(n416), .B(n415), .Z(n418) );
  XNOR2_X1 U470 ( .A(G29GAT), .B(G85GAT), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n418), .B(n417), .ZN(n419) );
  XNOR2_X1 U472 ( .A(n433), .B(n419), .ZN(n459) );
  XNOR2_X1 U473 ( .A(KEYINPUT91), .B(n459), .ZN(n506) );
  INV_X1 U474 ( .A(n506), .ZN(n558) );
  XOR2_X1 U475 ( .A(KEYINPUT22), .B(KEYINPUT88), .Z(n421) );
  XNOR2_X1 U476 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U478 ( .A(KEYINPUT87), .B(G162GAT), .Z(n423) );
  XNOR2_X1 U479 ( .A(G50GAT), .B(G22GAT), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n437) );
  XOR2_X1 U482 ( .A(G106GAT), .B(n426), .Z(n428) );
  NAND2_X1 U483 ( .A1(G228GAT), .A2(G233GAT), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U485 ( .A(n429), .B(G218GAT), .Z(n435) );
  XOR2_X1 U486 ( .A(G78GAT), .B(G148GAT), .Z(n431) );
  XNOR2_X1 U487 ( .A(KEYINPUT89), .B(KEYINPUT85), .ZN(n430) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U491 ( .A(n437), .B(n436), .ZN(n462) );
  AND2_X1 U492 ( .A1(n558), .A2(n462), .ZN(n438) );
  NAND2_X1 U493 ( .A1(n559), .A2(n438), .ZN(n440) );
  XOR2_X1 U494 ( .A(KEYINPUT118), .B(KEYINPUT55), .Z(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  NAND2_X1 U496 ( .A1(n553), .A2(n443), .ZN(n445) );
  NAND2_X1 U497 ( .A1(n553), .A2(n526), .ZN(n449) );
  XOR2_X1 U498 ( .A(KEYINPUT120), .B(KEYINPUT56), .Z(n447) );
  XNOR2_X1 U499 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n446) );
  XNOR2_X1 U500 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n449), .B(n448), .ZN(G1349GAT) );
  NAND2_X1 U502 ( .A1(n551), .A2(n450), .ZN(n484) );
  NOR2_X1 U503 ( .A1(n443), .A2(n544), .ZN(n451) );
  XNOR2_X1 U504 ( .A(n451), .B(KEYINPUT16), .ZN(n468) );
  INV_X1 U505 ( .A(n524), .ZN(n512) );
  NOR2_X1 U506 ( .A1(n462), .A2(n512), .ZN(n453) );
  XNOR2_X1 U507 ( .A(KEYINPUT26), .B(KEYINPUT96), .ZN(n452) );
  XNOR2_X1 U508 ( .A(n453), .B(n452), .ZN(n560) );
  XOR2_X1 U509 ( .A(KEYINPUT27), .B(n472), .Z(n461) );
  NAND2_X1 U510 ( .A1(n560), .A2(n461), .ZN(n458) );
  NOR2_X1 U511 ( .A1(n524), .A2(n472), .ZN(n454) );
  XNOR2_X1 U512 ( .A(KEYINPUT97), .B(n454), .ZN(n455) );
  NAND2_X1 U513 ( .A1(n455), .A2(n462), .ZN(n456) );
  XOR2_X1 U514 ( .A(KEYINPUT25), .B(n456), .Z(n457) );
  NAND2_X1 U515 ( .A1(n458), .A2(n457), .ZN(n460) );
  NAND2_X1 U516 ( .A1(n460), .A2(n459), .ZN(n467) );
  NAND2_X1 U517 ( .A1(n506), .A2(n461), .ZN(n520) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT64), .ZN(n463) );
  XNOR2_X1 U519 ( .A(n463), .B(KEYINPUT28), .ZN(n522) );
  NAND2_X1 U520 ( .A1(n524), .A2(n522), .ZN(n464) );
  NOR2_X1 U521 ( .A1(n520), .A2(n464), .ZN(n465) );
  XNOR2_X1 U522 ( .A(KEYINPUT95), .B(n465), .ZN(n466) );
  NAND2_X1 U523 ( .A1(n467), .A2(n466), .ZN(n478) );
  NAND2_X1 U524 ( .A1(n468), .A2(n478), .ZN(n495) );
  NOR2_X1 U525 ( .A1(n484), .A2(n495), .ZN(n469) );
  XNOR2_X1 U526 ( .A(KEYINPUT98), .B(n469), .ZN(n476) );
  NAND2_X1 U527 ( .A1(n476), .A2(n506), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n470), .B(KEYINPUT34), .ZN(n471) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n471), .ZN(G1324GAT) );
  INV_X1 U530 ( .A(n472), .ZN(n509) );
  NAND2_X1 U531 ( .A1(n476), .A2(n509), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n473), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U533 ( .A(G15GAT), .B(KEYINPUT35), .Z(n475) );
  NAND2_X1 U534 ( .A1(n476), .A2(n512), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(G1326GAT) );
  INV_X1 U536 ( .A(n522), .ZN(n515) );
  NAND2_X1 U537 ( .A1(n476), .A2(n515), .ZN(n477) );
  XNOR2_X1 U538 ( .A(n477), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U539 ( .A(G29GAT), .B(KEYINPUT39), .Z(n488) );
  XOR2_X1 U540 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n483) );
  NAND2_X1 U541 ( .A1(n544), .A2(n478), .ZN(n479) );
  XOR2_X1 U542 ( .A(KEYINPUT99), .B(n479), .Z(n480) );
  NOR2_X1 U543 ( .A1(n575), .A2(n480), .ZN(n481) );
  XNOR2_X1 U544 ( .A(n481), .B(KEYINPUT37), .ZN(n482) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n505) );
  NOR2_X1 U546 ( .A1(n505), .A2(n484), .ZN(n486) );
  XNOR2_X1 U547 ( .A(KEYINPUT102), .B(KEYINPUT38), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n493) );
  NAND2_X1 U549 ( .A1(n493), .A2(n506), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  XOR2_X1 U551 ( .A(G36GAT), .B(KEYINPUT103), .Z(n490) );
  NAND2_X1 U552 ( .A1(n493), .A2(n509), .ZN(n489) );
  XNOR2_X1 U553 ( .A(n490), .B(n489), .ZN(G1329GAT) );
  NAND2_X1 U554 ( .A1(n512), .A2(n493), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n491), .B(KEYINPUT40), .ZN(n492) );
  XNOR2_X1 U556 ( .A(G43GAT), .B(n492), .ZN(G1330GAT) );
  NAND2_X1 U557 ( .A1(n493), .A2(n515), .ZN(n494) );
  XNOR2_X1 U558 ( .A(G50GAT), .B(n494), .ZN(G1331GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT104), .B(KEYINPUT42), .Z(n497) );
  INV_X1 U560 ( .A(n563), .ZN(n537) );
  NAND2_X1 U561 ( .A1(n526), .A2(n537), .ZN(n504) );
  NOR2_X1 U562 ( .A1(n504), .A2(n495), .ZN(n501) );
  NAND2_X1 U563 ( .A1(n501), .A2(n506), .ZN(n496) );
  XNOR2_X1 U564 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U565 ( .A(G57GAT), .B(n498), .Z(G1332GAT) );
  NAND2_X1 U566 ( .A1(n501), .A2(n509), .ZN(n499) );
  XNOR2_X1 U567 ( .A(n499), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U568 ( .A1(n512), .A2(n501), .ZN(n500) );
  XNOR2_X1 U569 ( .A(n500), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U570 ( .A(G78GAT), .B(KEYINPUT43), .Z(n503) );
  NAND2_X1 U571 ( .A1(n501), .A2(n515), .ZN(n502) );
  XNOR2_X1 U572 ( .A(n503), .B(n502), .ZN(G1335GAT) );
  XOR2_X1 U573 ( .A(G85GAT), .B(KEYINPUT105), .Z(n508) );
  NOR2_X1 U574 ( .A1(n505), .A2(n504), .ZN(n516) );
  NAND2_X1 U575 ( .A1(n516), .A2(n506), .ZN(n507) );
  XNOR2_X1 U576 ( .A(n508), .B(n507), .ZN(G1336GAT) );
  NAND2_X1 U577 ( .A1(n516), .A2(n509), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n510), .B(KEYINPUT106), .ZN(n511) );
  XNOR2_X1 U579 ( .A(G92GAT), .B(n511), .ZN(G1337GAT) );
  XOR2_X1 U580 ( .A(G99GAT), .B(KEYINPUT107), .Z(n514) );
  NAND2_X1 U581 ( .A1(n516), .A2(n512), .ZN(n513) );
  XNOR2_X1 U582 ( .A(n514), .B(n513), .ZN(G1338GAT) );
  XOR2_X1 U583 ( .A(KEYINPUT108), .B(KEYINPUT44), .Z(n518) );
  NAND2_X1 U584 ( .A1(n516), .A2(n515), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(n519) );
  XOR2_X1 U586 ( .A(G106GAT), .B(n519), .Z(G1339GAT) );
  NOR2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n536) );
  NAND2_X1 U588 ( .A1(n522), .A2(n536), .ZN(n523) );
  NOR2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n533) );
  NAND2_X1 U590 ( .A1(n533), .A2(n551), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G113GAT), .B(n525), .ZN(G1340GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U593 ( .A1(n533), .A2(n526), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U595 ( .A(G120GAT), .B(n529), .Z(G1341GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT114), .B(KEYINPUT50), .Z(n531) );
  NAND2_X1 U597 ( .A1(n533), .A2(n570), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U599 ( .A(G127GAT), .B(n532), .Z(G1342GAT) );
  XOR2_X1 U600 ( .A(G134GAT), .B(KEYINPUT51), .Z(n535) );
  NAND2_X1 U601 ( .A1(n533), .A2(n443), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(G1343GAT) );
  NAND2_X1 U603 ( .A1(n560), .A2(n536), .ZN(n548) );
  NOR2_X1 U604 ( .A1(n537), .A2(n548), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G141GAT), .B(KEYINPUT115), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(G1344GAT) );
  NOR2_X1 U607 ( .A1(n540), .A2(n548), .ZN(n542) );
  XNOR2_X1 U608 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n541) );
  XNOR2_X1 U609 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(n543), .ZN(G1345GAT) );
  NOR2_X1 U611 ( .A1(n544), .A2(n548), .ZN(n546) );
  XNOR2_X1 U612 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n545) );
  XNOR2_X1 U613 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G155GAT), .B(n547), .ZN(G1346GAT) );
  NOR2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U616 ( .A(G162GAT), .B(n550), .Z(G1347GAT) );
  NAND2_X1 U617 ( .A1(n553), .A2(n551), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(n552), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(G183GAT), .B(KEYINPUT121), .Z(n555) );
  NAND2_X1 U620 ( .A1(n553), .A2(n570), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1350GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n557) );
  XNOR2_X1 U623 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n565) );
  AND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U627 ( .A(KEYINPUT122), .B(n562), .Z(n574) );
  NAND2_X1 U628 ( .A1(n574), .A2(n563), .ZN(n564) );
  XOR2_X1 U629 ( .A(n565), .B(n564), .Z(G1352GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT61), .B(KEYINPUT125), .Z(n567) );
  NAND2_X1 U631 ( .A1(n389), .A2(n574), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U633 ( .A(G204GAT), .B(KEYINPUT124), .Z(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1353GAT) );
  NAND2_X1 U635 ( .A1(n574), .A2(n570), .ZN(n571) );
  XNOR2_X1 U636 ( .A(n571), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n573) );
  XNOR2_X1 U638 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n572) );
  XNOR2_X1 U639 ( .A(n573), .B(n572), .ZN(n578) );
  INV_X1 U640 ( .A(n574), .ZN(n576) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(n578), .B(n577), .Z(G1355GAT) );
endmodule

