//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:28 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1247, new_n1248, new_n1249,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT0), .Z(new_n211));
  INV_X1    g0011(.A(G87), .ZN(new_n212));
  INV_X1    g0012(.A(G250), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G244), .ZN(new_n215));
  INV_X1    g0015(.A(G97), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  OAI22_X1  g0017(.A1(new_n202), .A2(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n214), .B(new_n218), .C1(G116), .C2(G270), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G50), .A2(G226), .ZN(new_n220));
  AND2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G58), .ZN(new_n222));
  INV_X1    g0022(.A(G232), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(G68), .ZN(new_n227));
  INV_X1    g0027(.A(G238), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n208), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n206), .ZN(new_n233));
  OAI21_X1  g0033(.A(G50), .B1(G58), .B2(G68), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(KEYINPUT64), .Z(new_n235));
  AOI211_X1 g0035(.A(new_n211), .B(new_n231), .C1(new_n233), .C2(new_n235), .ZN(G361));
  XOR2_X1   g0036(.A(G226), .B(G232), .Z(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G250), .B(G257), .Z(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G358));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XOR2_X1   g0046(.A(G50), .B(G58), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  OAI211_X1 g0052(.A(new_n205), .B(G274), .C1(G41), .C2(G45), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT66), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(KEYINPUT73), .ZN(new_n255));
  NAND2_X1  g0055(.A1(G33), .A2(G97), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT3), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n261), .B1(G232), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G226), .A2(G1698), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n256), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n232), .B1(G33), .B2(G41), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n265), .A2(new_n266), .B1(new_n270), .B2(G238), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n255), .A2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(KEYINPUT13), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT13), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n275), .B1(new_n255), .B2(new_n271), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G200), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(new_n232), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n206), .A2(new_n258), .A3(KEYINPUT67), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(G20), .B2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G50), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n258), .A2(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n290), .A2(new_n202), .B1(new_n206), .B2(G68), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n281), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT11), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n205), .A2(G13), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n206), .A2(G68), .ZN(new_n296));
  AOI21_X1  g0096(.A(KEYINPUT74), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  XOR2_X1   g0097(.A(new_n297), .B(KEYINPUT12), .Z(new_n298));
  AOI21_X1  g0098(.A(new_n281), .B1(new_n205), .B2(G20), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n298), .B1(G68), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n293), .A2(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n274), .A2(G190), .A3(new_n277), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n279), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(G169), .B1(new_n273), .B2(new_n276), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT14), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT14), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n308), .B(G169), .C1(new_n273), .C2(new_n276), .ZN(new_n309));
  INV_X1    g0109(.A(G179), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n307), .B(new_n309), .C1(new_n310), .C2(new_n278), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n305), .B1(new_n301), .B2(new_n311), .ZN(new_n312));
  XOR2_X1   g0112(.A(KEYINPUT8), .B(G58), .Z(new_n313));
  AOI22_X1  g0113(.A1(new_n289), .A2(new_n313), .B1(new_n285), .B2(G150), .ZN(new_n314));
  XNOR2_X1  g0114(.A(new_n314), .B(KEYINPUT68), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n201), .A2(new_n206), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n281), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n287), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n299), .A2(G50), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n317), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT9), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n270), .A2(G226), .ZN(new_n325));
  INV_X1    g0125(.A(new_n261), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n202), .ZN(new_n327));
  MUX2_X1   g0127(.A(G222), .B(G223), .S(G1698), .Z(new_n328));
  OAI211_X1 g0128(.A(new_n327), .B(new_n266), .C1(new_n326), .C2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n254), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n325), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G190), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(G200), .B2(new_n331), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n322), .A2(new_n323), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n324), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(KEYINPUT72), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT10), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n336), .B(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n331), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n322), .B1(G169), .B2(new_n341), .ZN(new_n342));
  OR2_X1    g0142(.A1(new_n342), .A2(KEYINPUT69), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(KEYINPUT69), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n343), .B(new_n344), .C1(G179), .C2(new_n331), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n318), .A2(G77), .ZN(new_n346));
  INV_X1    g0146(.A(new_n281), .ZN(new_n347));
  XOR2_X1   g0147(.A(KEYINPUT15), .B(G87), .Z(new_n348));
  AOI22_X1  g0148(.A1(new_n348), .A2(new_n289), .B1(G20), .B2(G77), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n313), .A2(new_n285), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n347), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AOI211_X1 g0151(.A(new_n346), .B(new_n351), .C1(G77), .C2(new_n299), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n228), .A2(G1698), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(G232), .B2(G1698), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n261), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT70), .B(G107), .ZN(new_n356));
  OAI211_X1 g0156(.A(new_n355), .B(new_n266), .C1(new_n261), .C2(new_n356), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n357), .B(new_n330), .C1(new_n215), .C2(new_n269), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G200), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n352), .B(new_n359), .C1(new_n332), .C2(new_n358), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n312), .A2(new_n340), .A3(new_n345), .A4(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n257), .A2(KEYINPUT75), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT75), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT3), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n364), .A3(G33), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n259), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(G226), .A3(G1698), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT77), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n258), .A2(new_n212), .ZN(new_n369));
  AOI21_X1  g0169(.A(G1698), .B1(new_n365), .B2(new_n259), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(G223), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT77), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n366), .A2(new_n372), .A3(G226), .A4(G1698), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n368), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n266), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n269), .A2(new_n223), .ZN(new_n376));
  INV_X1    g0176(.A(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n330), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(G200), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n375), .A2(G190), .A3(new_n330), .A4(new_n377), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n313), .A2(new_n319), .ZN(new_n381));
  INV_X1    g0181(.A(new_n299), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n381), .B1(new_n382), .B2(new_n313), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n222), .A2(new_n227), .ZN(new_n385));
  NOR2_X1   g0185(.A1(G58), .A2(G68), .ZN(new_n386));
  OAI21_X1  g0186(.A(G20), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(G159), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n387), .B1(new_n286), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT7), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n261), .B2(G20), .ZN(new_n391));
  XNOR2_X1  g0191(.A(KEYINPUT75), .B(KEYINPUT3), .ZN(new_n392));
  OAI211_X1 g0192(.A(KEYINPUT7), .B(new_n206), .C1(new_n392), .C2(G33), .ZN(new_n393));
  INV_X1    g0193(.A(new_n260), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n389), .B1(new_n395), .B2(G68), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT76), .B1(new_n396), .B2(KEYINPUT16), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n365), .A2(new_n206), .A3(new_n259), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n227), .B1(new_n398), .B2(KEYINPUT7), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n365), .A2(new_n390), .A3(new_n206), .A4(new_n259), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n389), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n347), .B1(new_n401), .B2(KEYINPUT16), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT76), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n362), .A2(new_n364), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n390), .B1(new_n405), .B2(new_n258), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n406), .A2(new_n206), .A3(new_n260), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n227), .B1(new_n407), .B2(new_n391), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n403), .B(new_n404), .C1(new_n408), .C2(new_n389), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n397), .A2(new_n402), .A3(new_n409), .ZN(new_n410));
  NAND4_X1  g0210(.A1(new_n379), .A2(new_n380), .A3(new_n384), .A4(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT17), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n384), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n415), .A2(KEYINPUT17), .A3(new_n380), .A4(new_n379), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n375), .A2(G179), .A3(new_n330), .A4(new_n377), .ZN(new_n417));
  AOI211_X1 g0217(.A(new_n254), .B(new_n376), .C1(new_n374), .C2(new_n266), .ZN(new_n418));
  INV_X1    g0218(.A(G169), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n420), .A2(new_n414), .A3(KEYINPUT18), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(KEYINPUT18), .B1(new_n420), .B2(new_n414), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n413), .B(new_n416), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n358), .A2(G179), .ZN(new_n425));
  XOR2_X1   g0225(.A(new_n425), .B(KEYINPUT71), .Z(new_n426));
  INV_X1    g0226(.A(new_n352), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n358), .A2(new_n419), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NOR3_X1   g0230(.A1(new_n361), .A2(new_n424), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n205), .A2(G33), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n318), .A2(new_n432), .A3(new_n232), .A4(new_n280), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(KEYINPUT82), .A3(G116), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT82), .ZN(new_n436));
  INV_X1    g0236(.A(G116), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n436), .B1(new_n433), .B2(new_n437), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n280), .A2(new_n232), .B1(G20), .B2(new_n437), .ZN(new_n440));
  NAND2_X1  g0240(.A1(G33), .A2(G283), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(new_n206), .C1(G33), .C2(new_n216), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(KEYINPUT20), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(KEYINPUT20), .B1(new_n440), .B2(new_n442), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n437), .A2(G20), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n444), .A2(new_n445), .B1(new_n294), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(G179), .B1(new_n439), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(G41), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n449), .A2(KEYINPUT5), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT5), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n205), .B(G45), .C1(new_n451), .C2(G41), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n267), .B(G270), .C1(new_n450), .C2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n450), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G274), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n365), .A2(new_n259), .B1(new_n217), .B2(new_n262), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n225), .A2(G1698), .ZN(new_n457));
  AOI22_X1  g0257(.A1(new_n456), .A2(new_n457), .B1(G303), .B2(new_n326), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n453), .B(new_n455), .C1(new_n458), .C2(new_n267), .ZN(new_n459));
  OAI21_X1  g0259(.A(KEYINPUT83), .B1(new_n448), .B2(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n217), .A2(new_n262), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n366), .A2(new_n461), .A3(new_n457), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n326), .A2(G303), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n267), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(new_n453), .ZN(new_n465));
  INV_X1    g0265(.A(new_n455), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n294), .A2(new_n446), .ZN(new_n468));
  INV_X1    g0268(.A(new_n445), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n468), .B1(new_n469), .B2(new_n443), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n435), .A2(new_n438), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n310), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT83), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n467), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n470), .A2(new_n471), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n459), .A2(new_n475), .A3(KEYINPUT21), .A4(G169), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n460), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(KEYINPUT84), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT21), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n475), .A2(G169), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n479), .B1(new_n480), .B2(new_n467), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT84), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n460), .A2(new_n474), .A3(new_n482), .A4(new_n476), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n459), .A2(G200), .ZN(new_n484));
  INV_X1    g0284(.A(new_n475), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n484), .B(new_n485), .C1(new_n332), .C2(new_n459), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n478), .A2(new_n481), .A3(new_n483), .A4(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT24), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n212), .A2(G20), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n261), .A2(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT22), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI21_X1  g0292(.A(KEYINPUT23), .B1(new_n356), .B2(new_n206), .ZN(new_n493));
  NOR3_X1   g0293(.A1(new_n258), .A2(new_n437), .A3(G20), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n206), .A2(KEYINPUT23), .A3(G107), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n492), .A2(new_n493), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n366), .A2(KEYINPUT22), .A3(new_n489), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n488), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AOI211_X1 g0300(.A(new_n494), .B(new_n496), .C1(new_n490), .C2(new_n491), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n366), .A2(KEYINPUT22), .A3(new_n489), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n501), .A2(KEYINPUT24), .A3(new_n493), .A4(new_n502), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n500), .A2(new_n503), .A3(new_n281), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n434), .A2(G107), .ZN(new_n505));
  AND2_X1   g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n454), .A2(new_n266), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G264), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n365), .A2(new_n259), .B1(new_n213), .B2(new_n262), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n217), .A2(G1698), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n509), .A2(new_n510), .B1(G33), .B2(G294), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n455), .B(new_n508), .C1(new_n511), .C2(new_n267), .ZN(new_n512));
  OR2_X1    g0312(.A1(new_n512), .A2(new_n332), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n318), .A2(G107), .ZN(new_n514));
  XNOR2_X1  g0314(.A(KEYINPUT85), .B(KEYINPUT25), .ZN(new_n515));
  XNOR2_X1  g0315(.A(new_n514), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n512), .A2(G200), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n506), .A2(new_n513), .A3(new_n516), .A4(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n262), .A2(KEYINPUT4), .A3(G244), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(new_n213), .B2(new_n262), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n261), .ZN(new_n521));
  AOI211_X1 g0321(.A(new_n215), .B(G1698), .C1(new_n365), .C2(new_n259), .ZN(new_n522));
  XOR2_X1   g0322(.A(KEYINPUT79), .B(KEYINPUT4), .Z(new_n523));
  OAI211_X1 g0323(.A(new_n441), .B(new_n521), .C1(new_n522), .C2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(new_n266), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n267), .B1(new_n450), .B2(new_n452), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n455), .B1(new_n526), .B2(new_n217), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n419), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n318), .A2(new_n216), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(new_n434), .B2(new_n216), .ZN(new_n532));
  XNOR2_X1  g0332(.A(new_n532), .B(KEYINPUT78), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n286), .A2(new_n202), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n224), .A2(KEYINPUT6), .A3(G97), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n216), .A2(new_n224), .ZN(new_n536));
  NOR2_X1   g0336(.A1(G97), .A2(G107), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n535), .B1(new_n538), .B2(KEYINPUT6), .ZN(new_n539));
  AOI221_X4 g0339(.A(new_n534), .B1(G20), .B2(new_n539), .C1(new_n395), .C2(new_n356), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n533), .B1(new_n540), .B2(new_n347), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n527), .B1(new_n524), .B2(new_n266), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n310), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n530), .A2(new_n541), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n529), .A2(G200), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT78), .ZN(new_n546));
  XNOR2_X1  g0346(.A(new_n532), .B(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n395), .A2(new_n356), .B1(G20), .B2(new_n539), .ZN(new_n548));
  INV_X1    g0348(.A(new_n534), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n547), .B1(new_n550), .B2(new_n281), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n542), .A2(G190), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n545), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n504), .A2(new_n505), .A3(new_n516), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n512), .A2(new_n419), .ZN(new_n555));
  OR2_X1    g0355(.A1(new_n512), .A2(G179), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n518), .A2(new_n544), .A3(new_n553), .A4(new_n557), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n205), .A2(G45), .A3(G274), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(G45), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n267), .B(G250), .C1(G1), .C2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n258), .A2(new_n437), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n262), .A2(G244), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n564), .B1(new_n365), .B2(new_n259), .ZN(new_n565));
  NOR2_X1   g0365(.A1(G238), .A2(G1698), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n563), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n560), .B(new_n562), .C1(new_n568), .C2(new_n267), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G169), .ZN(new_n570));
  AOI211_X1 g0370(.A(new_n566), .B(new_n564), .C1(new_n365), .C2(new_n259), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n266), .B1(new_n571), .B2(new_n563), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n572), .A2(G179), .A3(new_n560), .A4(new_n562), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(KEYINPUT80), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n366), .A2(new_n206), .A3(G68), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT19), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n577), .B1(new_n290), .B2(new_n216), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n206), .B1(new_n256), .B2(new_n577), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n212), .A2(new_n216), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n579), .B1(new_n356), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n576), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT81), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n576), .A2(KEYINPUT81), .A3(new_n578), .A4(new_n581), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n584), .A2(new_n281), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n348), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n319), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n434), .A2(new_n348), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT80), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n570), .A2(new_n591), .A3(new_n573), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n575), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  AND2_X1   g0393(.A1(new_n586), .A2(new_n588), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n569), .A2(new_n332), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n569), .A2(G200), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n434), .A2(G87), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n594), .A2(new_n596), .A3(new_n597), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n593), .A2(new_n599), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n487), .A2(new_n558), .A3(new_n600), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n431), .A2(new_n601), .ZN(G372));
  NAND3_X1  g0402(.A1(new_n518), .A2(new_n544), .A3(new_n553), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n590), .A2(new_n574), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n586), .A2(new_n597), .A3(new_n598), .A4(new_n588), .ZN(new_n605));
  OAI21_X1  g0405(.A(new_n604), .B1(new_n595), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT86), .B1(new_n603), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(new_n557), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n481), .A2(new_n460), .A3(new_n476), .A4(new_n474), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AND2_X1   g0410(.A1(new_n553), .A2(new_n544), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT86), .ZN(new_n612));
  AND4_X1   g0412(.A1(new_n597), .A2(new_n586), .A3(new_n598), .A4(new_n588), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n613), .A2(new_n596), .B1(new_n574), .B2(new_n590), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n611), .A2(new_n612), .A3(new_n518), .A4(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n607), .A2(new_n610), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n604), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT26), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n606), .B2(new_n544), .ZN(new_n619));
  AOI21_X1  g0419(.A(G169), .B1(new_n525), .B2(new_n528), .ZN(new_n620));
  AOI211_X1 g0420(.A(G179), .B(new_n527), .C1(new_n524), .C2(new_n266), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n551), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  XOR2_X1   g0422(.A(KEYINPUT87), .B(KEYINPUT26), .Z(new_n623));
  NAND4_X1  g0423(.A1(new_n593), .A2(new_n599), .A3(new_n622), .A4(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n617), .B1(new_n619), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n616), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n431), .A2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(new_n345), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n311), .A2(new_n301), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n429), .ZN(new_n630));
  XNOR2_X1  g0430(.A(new_n411), .B(KEYINPUT17), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(new_n631), .A3(new_n304), .ZN(new_n632));
  INV_X1    g0432(.A(new_n423), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n421), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n628), .B1(new_n635), .B2(new_n340), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n627), .A2(new_n636), .ZN(G369));
  NAND2_X1  g0437(.A1(new_n295), .A2(new_n206), .ZN(new_n638));
  OR3_X1    g0438(.A1(new_n638), .A2(KEYINPUT88), .A3(KEYINPUT27), .ZN(new_n639));
  INV_X1    g0439(.A(G213), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n640), .B1(new_n638), .B2(KEYINPUT27), .ZN(new_n641));
  OAI21_X1  g0441(.A(KEYINPUT88), .B1(new_n638), .B2(KEYINPUT27), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n639), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(G343), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n475), .ZN(new_n646));
  XOR2_X1   g0446(.A(new_n646), .B(KEYINPUT89), .Z(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n609), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n487), .B2(new_n647), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(KEYINPUT90), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT90), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n648), .B(new_n651), .C1(new_n487), .C2(new_n647), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  AND4_X1   g0453(.A1(new_n505), .A2(new_n517), .A3(new_n504), .A4(new_n516), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n654), .A2(new_n513), .B1(new_n554), .B2(new_n645), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n655), .A2(new_n608), .ZN(new_n656));
  INV_X1    g0456(.A(new_n645), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n608), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n653), .A2(G330), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n478), .A2(new_n481), .A3(new_n483), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n662), .A2(new_n557), .A3(new_n657), .A4(new_n655), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(new_n658), .A3(new_n663), .ZN(G399));
  INV_X1    g0464(.A(new_n209), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n665), .A2(G41), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n356), .A2(G116), .A3(new_n580), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g0468(.A1(new_n666), .A2(new_n205), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT91), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n669), .A2(new_n670), .ZN(new_n672));
  INV_X1    g0472(.A(new_n666), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n671), .B(new_n672), .C1(new_n234), .C2(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT28), .ZN(new_n675));
  AOI211_X1 g0475(.A(KEYINPUT29), .B(new_n645), .C1(new_n616), .C2(new_n625), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT92), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n606), .A2(new_n544), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n593), .A2(new_n599), .A3(new_n622), .ZN(new_n679));
  INV_X1    g0479(.A(new_n623), .ZN(new_n680));
  AOI22_X1  g0480(.A1(new_n678), .A2(KEYINPUT26), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n677), .B1(new_n681), .B2(new_n617), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n606), .A2(new_n618), .A3(new_n544), .ZN(new_n684));
  OAI211_X1 g0484(.A(KEYINPUT92), .B(new_n604), .C1(new_n683), .C2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n603), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n686), .B(new_n614), .C1(new_n662), .C2(new_n608), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n682), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n657), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n676), .B1(new_n689), .B2(KEYINPUT29), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n558), .A2(new_n600), .ZN(new_n691));
  INV_X1    g0491(.A(new_n487), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n691), .A2(new_n692), .A3(new_n657), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT30), .ZN(new_n694));
  OR2_X1    g0494(.A1(new_n573), .A2(new_n459), .ZN(new_n695));
  INV_X1    g0495(.A(new_n511), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n696), .A2(new_n266), .B1(G264), .B2(new_n507), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n542), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n694), .B1(new_n695), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n573), .A2(new_n459), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n542), .A3(KEYINPUT30), .A4(new_n697), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n542), .A2(new_n467), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n702), .A2(new_n310), .A3(new_n569), .A4(new_n512), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n699), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n645), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT31), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(KEYINPUT31), .A3(new_n645), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n693), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(G330), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n690), .A2(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n675), .B1(new_n712), .B2(G1), .ZN(G364));
  NOR2_X1   g0513(.A1(G13), .A2(G33), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G20), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n232), .B1(G20), .B2(new_n419), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n665), .A2(new_n366), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n719), .B1(new_n561), .B2(new_n235), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n248), .A2(G45), .ZN(new_n721));
  AOI22_X1  g0521(.A1(new_n720), .A2(new_n721), .B1(new_n437), .B2(new_n665), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n209), .A2(new_n261), .ZN(new_n723));
  XOR2_X1   g0523(.A(new_n723), .B(KEYINPUT93), .Z(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G355), .ZN(new_n725));
  AOI211_X1 g0525(.A(new_n716), .B(new_n717), .C1(new_n722), .C2(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(G13), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n205), .B1(new_n728), .B2(G45), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n666), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n206), .A2(G190), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n310), .A2(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G200), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n310), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n733), .ZN(new_n738));
  OAI221_X1 g0538(.A(new_n261), .B1(new_n735), .B2(new_n202), .C1(new_n227), .C2(new_n738), .ZN(new_n739));
  NOR4_X1   g0539(.A1(new_n206), .A2(G179), .A3(G190), .A4(G200), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n740), .A2(KEYINPUT95), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(KEYINPUT95), .ZN(new_n742));
  AND2_X1   g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G159), .ZN(new_n744));
  XOR2_X1   g0544(.A(new_n744), .B(KEYINPUT32), .Z(new_n745));
  NOR2_X1   g0545(.A1(new_n736), .A2(G179), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(new_n733), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT96), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(G107), .ZN(new_n750));
  NOR3_X1   g0550(.A1(new_n332), .A2(G179), .A3(G200), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n206), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G97), .ZN(new_n754));
  NAND2_X1  g0554(.A1(G20), .A2(G190), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n734), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g0557(.A(new_n757), .B(KEYINPUT94), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n746), .A2(new_n756), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI22_X1  g0561(.A1(new_n759), .A2(G58), .B1(G87), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g0562(.A1(new_n745), .A2(new_n750), .A3(new_n754), .A4(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n737), .A2(new_n756), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n739), .B(new_n763), .C1(G50), .C2(new_n765), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT97), .Z(new_n767));
  INV_X1    g0567(.A(G326), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n764), .A2(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G283), .A2(new_n749), .B1(new_n743), .B2(G329), .ZN(new_n770));
  XOR2_X1   g0570(.A(new_n760), .B(KEYINPUT98), .Z(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G303), .ZN(new_n773));
  INV_X1    g0573(.A(G311), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n326), .B1(new_n735), .B2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G294), .ZN(new_n776));
  INV_X1    g0576(.A(G322), .ZN(new_n777));
  OAI22_X1  g0577(.A1(new_n752), .A2(new_n776), .B1(new_n757), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n738), .ZN(new_n779));
  XNOR2_X1  g0579(.A(KEYINPUT33), .B(G317), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n775), .B(new_n778), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n770), .A2(new_n773), .A3(new_n781), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n767), .B1(new_n769), .B2(new_n782), .ZN(new_n783));
  AOI211_X1 g0583(.A(new_n726), .B(new_n732), .C1(new_n783), .C2(new_n717), .ZN(new_n784));
  INV_X1    g0584(.A(new_n716), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n649), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n650), .A2(G330), .A3(new_n652), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(new_n732), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n653), .A2(G330), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n786), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT99), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(G396));
  AOI21_X1  g0592(.A(new_n645), .B1(new_n616), .B2(new_n625), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n360), .B1(new_n352), .B2(new_n657), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n429), .A2(new_n794), .ZN(new_n795));
  NAND4_X1  g0595(.A1(new_n426), .A2(new_n427), .A3(new_n428), .A4(new_n657), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  AOI211_X1 g0599(.A(new_n645), .B(new_n797), .C1(new_n616), .C2(new_n625), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(new_n710), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n732), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n797), .A2(new_n714), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n779), .A2(G150), .B1(new_n765), .B2(G137), .ZN(new_n805));
  INV_X1    g0605(.A(G143), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n805), .B1(new_n388), .B2(new_n735), .C1(new_n806), .C2(new_n758), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT34), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n749), .A2(G68), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n772), .A2(G50), .B1(new_n743), .B2(G132), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n808), .A2(new_n366), .A3(new_n809), .A4(new_n810), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n752), .A2(new_n222), .ZN(new_n812));
  INV_X1    g0612(.A(G283), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n754), .B1(new_n437), .B2(new_n735), .C1(new_n813), .C2(new_n738), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n261), .B(new_n814), .C1(G303), .C2(new_n765), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n772), .A2(G107), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n748), .A2(new_n212), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(new_n743), .B2(G311), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n815), .A2(new_n816), .A3(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n757), .A2(new_n776), .ZN(new_n820));
  OAI22_X1  g0620(.A1(new_n811), .A2(new_n812), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n717), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n717), .A2(new_n714), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n202), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n804), .A2(new_n731), .A3(new_n822), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n803), .A2(new_n825), .ZN(G384));
  INV_X1    g0626(.A(KEYINPUT38), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n401), .A2(KEYINPUT16), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(new_n281), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n401), .A2(KEYINPUT16), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n384), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT100), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI211_X1 g0633(.A(KEYINPUT100), .B(new_n384), .C1(new_n829), .C2(new_n830), .ZN(new_n834));
  AND2_X1   g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n643), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n631), .B2(new_n634), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n420), .A2(new_n414), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n414), .A2(new_n836), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT37), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n839), .A2(new_n411), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n417), .B(new_n643), .C1(new_n418), .C2(new_n419), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n833), .A2(new_n844), .A3(new_n834), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n841), .B1(new_n845), .B2(new_n411), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n827), .B1(new_n838), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n837), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n424), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n845), .A2(new_n411), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n842), .B1(new_n851), .B2(new_n841), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n850), .A2(new_n852), .A3(KEYINPUT38), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n848), .A2(KEYINPUT101), .A3(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT101), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n855), .B(new_n827), .C1(new_n838), .C2(new_n847), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT40), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n301), .A2(new_n645), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n629), .A2(new_n304), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n311), .A2(new_n301), .A3(new_n645), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n797), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n707), .A2(KEYINPUT102), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT102), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n705), .A2(new_n864), .A3(new_n706), .ZN(new_n865));
  NAND4_X1  g0665(.A1(new_n693), .A2(new_n863), .A3(new_n708), .A4(new_n865), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n862), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n857), .A2(new_n858), .A3(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n840), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n839), .A2(new_n411), .A3(new_n840), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT37), .ZN(new_n871));
  AOI22_X1  g0671(.A1(new_n424), .A2(new_n869), .B1(new_n842), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n853), .B1(new_n872), .B2(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n867), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(KEYINPUT40), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n876), .A2(new_n866), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(G330), .ZN(new_n878));
  INV_X1    g0678(.A(G330), .ZN(new_n879));
  INV_X1    g0679(.A(new_n708), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n601), .B2(new_n657), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n864), .B1(new_n705), .B2(new_n706), .ZN(new_n882));
  AOI211_X1 g0682(.A(KEYINPUT102), .B(KEYINPUT31), .C1(new_n704), .C2(new_n645), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n879), .B1(new_n881), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n431), .A2(new_n885), .ZN(new_n886));
  AOI22_X1  g0686(.A1(new_n877), .A2(new_n431), .B1(new_n878), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n854), .A2(KEYINPUT39), .A3(new_n856), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT39), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n853), .B(new_n889), .C1(KEYINPUT38), .C2(new_n872), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n629), .A2(new_n645), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n634), .A2(new_n836), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n860), .A2(new_n861), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n793), .A2(new_n798), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n896), .B1(new_n897), .B2(new_n796), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n894), .B1(new_n857), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g0700(.A(new_n887), .B(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT29), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n902), .B1(new_n688), .B2(new_n657), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n431), .B1(new_n903), .B2(new_n676), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n636), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n901), .B(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n205), .B2(new_n728), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n437), .B1(new_n539), .B2(KEYINPUT35), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n908), .B(new_n233), .C1(KEYINPUT35), .C2(new_n539), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n909), .B(KEYINPUT36), .ZN(new_n910));
  OAI21_X1  g0710(.A(G77), .B1(new_n222), .B2(new_n227), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n911), .A2(new_n234), .B1(G50), .B2(new_n227), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n912), .A2(G1), .A3(new_n727), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n907), .A2(new_n910), .A3(new_n913), .ZN(G367));
  NAND2_X1  g0714(.A1(new_n622), .A2(new_n657), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n541), .A2(new_n645), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n553), .A2(new_n544), .A3(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT42), .B1(new_n663), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n663), .A2(new_n658), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n658), .A2(KEYINPUT42), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n915), .B(new_n918), .C1(new_n921), .C2(new_n917), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n594), .A2(new_n598), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n645), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n614), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n604), .B2(new_n924), .ZN(new_n926));
  OR2_X1    g0726(.A1(new_n926), .A2(KEYINPUT43), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(KEYINPUT43), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n922), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT104), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n929), .B(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n922), .A2(new_n927), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT103), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n622), .A2(new_n645), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n917), .A2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n661), .A2(new_n937), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n934), .B(new_n938), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n666), .B(KEYINPUT41), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n919), .A2(new_n937), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT44), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n919), .A2(KEYINPUT44), .A3(new_n937), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n663), .A2(new_n658), .A3(new_n936), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT45), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n663), .A2(KEYINPUT45), .A3(new_n658), .A4(new_n936), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n944), .A2(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n950), .A2(KEYINPUT105), .A3(new_n661), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n787), .A2(new_n659), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n948), .A2(new_n949), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT44), .B1(new_n919), .B2(new_n937), .ZN(new_n954));
  AOI211_X1 g0754(.A(new_n943), .B(new_n936), .C1(new_n663), .C2(new_n658), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT105), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n952), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n951), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT106), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n663), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n787), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n660), .B1(new_n662), .B2(new_n657), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n650), .A2(new_n961), .A3(G330), .A4(new_n652), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n963), .B2(new_n965), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT107), .ZN(new_n969));
  NAND4_X1  g0769(.A1(new_n959), .A2(new_n712), .A3(new_n968), .A4(new_n969), .ZN(new_n970));
  OAI211_X1 g0770(.A(new_n690), .B(new_n710), .C1(new_n966), .C2(new_n967), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n661), .B1(new_n950), .B2(KEYINPUT105), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n956), .A2(new_n957), .A3(new_n952), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(KEYINPUT107), .B1(new_n971), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n941), .B1(new_n976), .B2(new_n712), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n939), .B1(new_n977), .B2(new_n730), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n752), .A2(new_n227), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(G150), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n980), .B1(new_n202), .B2(new_n747), .C1(new_n981), .C2(new_n757), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n326), .B1(new_n743), .B2(G137), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n806), .B2(new_n764), .ZN(new_n984));
  AOI211_X1 g0784(.A(new_n982), .B(new_n984), .C1(G58), .C2(new_n761), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n985), .B1(new_n287), .B2(new_n735), .C1(new_n388), .C2(new_n738), .ZN(new_n986));
  OAI21_X1  g0786(.A(KEYINPUT46), .B1(new_n771), .B2(new_n437), .ZN(new_n987));
  OR3_X1    g0787(.A1(new_n760), .A2(KEYINPUT46), .A3(new_n437), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n987), .A2(new_n988), .B1(new_n356), .B2(new_n753), .ZN(new_n989));
  INV_X1    g0789(.A(G303), .ZN(new_n990));
  INV_X1    g0790(.A(G317), .ZN(new_n991));
  INV_X1    g0791(.A(new_n743), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n989), .B1(new_n990), .B2(new_n758), .C1(new_n991), .C2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n735), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n993), .B1(G283), .B2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n747), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n366), .B1(G97), .B2(new_n996), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n995), .B(new_n997), .C1(new_n774), .C2(new_n764), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n738), .A2(new_n776), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n986), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT47), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n717), .ZN(new_n1002));
  OR2_X1    g0802(.A1(new_n926), .A2(new_n785), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n716), .A2(new_n717), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n209), .B2(new_n587), .C1(new_n719), .C2(new_n244), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1002), .A2(new_n731), .A3(new_n1003), .A4(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n978), .A2(new_n1006), .ZN(G387));
  NAND2_X1  g0807(.A1(new_n313), .A2(new_n287), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT50), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n667), .B1(new_n227), .B2(new_n202), .ZN(new_n1010));
  NOR3_X1   g0810(.A1(new_n1009), .A2(G45), .A3(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n718), .B1(new_n241), .B2(new_n561), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n724), .A2(new_n668), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n209), .A2(G107), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1004), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n731), .B(new_n1016), .C1(new_n660), .C2(new_n785), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n992), .A2(new_n981), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n764), .A2(new_n388), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n760), .A2(new_n202), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n313), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1021), .A2(new_n738), .B1(new_n287), .B2(new_n757), .ZN(new_n1022));
  NOR4_X1   g0822(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n753), .A2(new_n348), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n749), .A2(G97), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n366), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G68), .B2(new_n994), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1023), .A2(new_n1024), .A3(new_n1025), .A4(new_n1027), .ZN(new_n1028));
  AOI22_X1  g0828(.A1(G311), .A2(new_n779), .B1(new_n994), .B2(G303), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n777), .B2(new_n764), .C1(new_n758), .C2(new_n991), .ZN(new_n1030));
  XOR2_X1   g0830(.A(KEYINPUT108), .B(KEYINPUT48), .Z(new_n1031));
  XNOR2_X1  g0831(.A(new_n1030), .B(new_n1031), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n813), .B2(new_n752), .C1(new_n776), .C2(new_n760), .ZN(new_n1033));
  XOR2_X1   g0833(.A(new_n1033), .B(KEYINPUT49), .Z(new_n1034));
  OAI221_X1 g0834(.A(new_n1026), .B1(new_n437), .B2(new_n747), .C1(new_n992), .C2(new_n768), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1028), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT109), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1017), .B1(new_n1037), .B2(new_n717), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n968), .B2(new_n730), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n666), .B1(new_n712), .B2(new_n968), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n971), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(G393));
  INV_X1    g0842(.A(KEYINPUT110), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n661), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n952), .A2(KEYINPUT110), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1044), .A2(new_n950), .A3(new_n1045), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n956), .A2(new_n1043), .A3(new_n661), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(KEYINPUT111), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT111), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1046), .A2(new_n1050), .A3(new_n1047), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n730), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n732), .B1(new_n937), .B2(new_n716), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G107), .A2(new_n749), .B1(new_n743), .B2(G322), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n752), .A2(new_n437), .B1(new_n735), .B2(new_n776), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n261), .B(new_n1055), .C1(G303), .C2(new_n779), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n761), .A2(G283), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n764), .A2(new_n991), .B1(new_n757), .B2(new_n774), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT52), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1054), .A2(new_n1056), .A3(new_n1057), .A4(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n764), .A2(new_n981), .B1(new_n757), .B2(new_n388), .ZN(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT113), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n1062), .B(KEYINPUT51), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n817), .B1(new_n743), .B2(G143), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n753), .A2(G77), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n287), .B2(new_n738), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1026), .B(new_n1066), .C1(G68), .C2(new_n761), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1063), .A2(new_n1064), .A3(new_n1067), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n1021), .A2(new_n735), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1060), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n717), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1004), .B1(new_n216), .B2(new_n209), .C1(new_n719), .C2(new_n251), .ZN(new_n1072));
  XOR2_X1   g0872(.A(new_n1072), .B(KEYINPUT112), .Z(new_n1073));
  NAND3_X1  g0873(.A1(new_n1053), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1052), .A2(new_n1074), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1041), .A2(new_n1048), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n970), .B2(new_n975), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1075), .B1(new_n1077), .B2(new_n666), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(G390));
  AND3_X1   g0879(.A1(new_n862), .A2(new_n866), .A3(G330), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n888), .B(new_n890), .C1(new_n898), .C2(new_n892), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n688), .A2(new_n657), .A3(new_n795), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n896), .B1(new_n1083), .B2(new_n796), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n892), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n873), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1080), .B1(new_n1082), .B2(new_n1087), .ZN(new_n1088));
  OR2_X1    g0888(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n862), .A2(G330), .A3(new_n709), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1089), .A2(new_n1081), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1088), .A2(new_n730), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n888), .A2(new_n714), .A3(new_n890), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1065), .B1(new_n437), .B2(new_n757), .C1(new_n813), .C2(new_n764), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n261), .B(new_n1094), .C1(G97), .C2(new_n994), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n779), .A2(new_n356), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n772), .A2(G87), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(G68), .A2(new_n749), .B1(new_n743), .B2(G294), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(G125), .ZN(new_n1100));
  OAI221_X1 g0900(.A(new_n261), .B1(new_n287), .B2(new_n747), .C1(new_n992), .C2(new_n1100), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT117), .Z(new_n1102));
  XOR2_X1   g0902(.A(KEYINPUT54), .B(G143), .Z(new_n1103));
  AOI22_X1  g0903(.A1(G137), .A2(new_n779), .B1(new_n994), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT115), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1106), .B(new_n1107), .C1(new_n388), .C2(new_n752), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT116), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n760), .A2(new_n981), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT53), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1102), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g0912(.A(G128), .ZN(new_n1113));
  INV_X1    g0913(.A(G132), .ZN(new_n1114));
  OAI22_X1  g0914(.A1(new_n764), .A2(new_n1113), .B1(new_n757), .B2(new_n1114), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT118), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1099), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n717), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n823), .A2(new_n1021), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1093), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1092), .B1(new_n732), .B2(new_n1120), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1089), .A2(new_n1081), .A3(new_n1090), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n885), .A2(new_n862), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n1089), .B2(new_n1081), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n796), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1126), .B1(new_n793), .B2(new_n798), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n896), .B1(new_n710), .B2(new_n797), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1127), .B1(new_n1128), .B2(new_n1123), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT114), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n798), .B1(new_n885), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n866), .A2(G330), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1132), .A2(KEYINPUT114), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n896), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1083), .A2(new_n796), .A3(new_n1090), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1129), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n904), .A2(new_n636), .A3(new_n886), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n673), .B1(new_n1125), .B2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1128), .A2(new_n1123), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n897), .A2(new_n796), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n797), .B1(new_n1132), .B2(KEYINPUT114), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n885), .A2(new_n1130), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n895), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1143), .B1(new_n1146), .B2(new_n1135), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n904), .A2(new_n636), .A3(new_n886), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1121), .B1(new_n1140), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(G378));
  INV_X1    g0952(.A(KEYINPUT121), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n340), .A2(new_n345), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n322), .A2(new_n836), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n340), .A2(new_n345), .A3(new_n1155), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1159), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n893), .A2(new_n899), .A3(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n879), .B1(new_n868), .B2(new_n875), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1085), .B1(new_n888), .B2(new_n890), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n894), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n854), .A2(new_n856), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n895), .B1(new_n800), .B2(new_n1126), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1162), .B1(new_n1166), .B2(new_n1170), .ZN(new_n1171));
  AND3_X1   g0971(.A1(new_n1164), .A2(new_n1165), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1165), .B1(new_n1164), .B2(new_n1171), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1153), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1088), .A2(new_n1139), .A3(new_n1091), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n1148), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1163), .B1(new_n893), .B2(new_n899), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1166), .A2(new_n1170), .A3(new_n1162), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n878), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1164), .A2(new_n1165), .A3(new_n1171), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(KEYINPUT121), .A3(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1174), .A2(new_n1176), .A3(new_n1181), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT57), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1176), .B(KEYINPUT57), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1184), .A2(new_n666), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT122), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1174), .A2(new_n730), .A3(new_n1181), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1162), .A2(new_n714), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n752), .A2(new_n981), .B1(new_n764), .B2(new_n1100), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(G132), .A2(new_n779), .B1(new_n994), .B2(G137), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n1113), .B2(new_n757), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1190), .B(new_n1192), .C1(new_n761), .C2(new_n1103), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1194));
  XNOR2_X1  g0994(.A(new_n1193), .B(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(KEYINPUT120), .B(G124), .ZN(new_n1196));
  AOI21_X1  g0996(.A(G41), .B1(new_n743), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(G33), .B1(new_n996), .B2(G159), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1195), .A2(new_n1197), .A3(new_n1198), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n366), .B(new_n1020), .C1(new_n743), .C2(G283), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n587), .A2(new_n735), .B1(new_n216), .B2(new_n738), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n449), .B1(new_n757), .B2(new_n224), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n747), .A2(new_n222), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n764), .A2(new_n437), .ZN(new_n1204));
  NOR4_X1   g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1200), .A2(new_n980), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT58), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(G41), .B1(new_n392), .B2(G33), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1199), .B(new_n1208), .C1(G50), .C2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n717), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n823), .A2(new_n287), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1189), .A2(new_n731), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1187), .B1(new_n1188), .B2(new_n1214), .ZN(new_n1215));
  AND3_X1   g1015(.A1(new_n1188), .A2(new_n1187), .A3(new_n1214), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1186), .B1(new_n1215), .B2(new_n1216), .ZN(G375));
  NAND2_X1  g1017(.A1(new_n896), .A2(new_n714), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n772), .A2(G97), .B1(new_n749), .B2(G77), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1219), .B1(new_n992), .B2(new_n990), .ZN(new_n1220));
  OAI221_X1 g1020(.A(new_n1024), .B1(new_n437), .B2(new_n738), .C1(new_n813), .C2(new_n757), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1222), .B(new_n326), .C1(new_n776), .C2(new_n764), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1220), .B(new_n1223), .C1(new_n356), .C2(new_n994), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n759), .A2(G137), .B1(G132), .B2(new_n765), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n388), .B2(new_n771), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1203), .B1(new_n743), .B2(G128), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1026), .B1(new_n779), .B2(new_n1103), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(new_n981), .C2(new_n735), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1226), .B(new_n1229), .C1(G50), .C2(new_n753), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n717), .B1(new_n1224), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n823), .A2(new_n227), .ZN(new_n1232));
  AND4_X1   g1032(.A1(new_n731), .A2(new_n1218), .A3(new_n1231), .A4(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1233), .B1(new_n1147), .B2(new_n730), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n940), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1234), .B1(new_n1235), .B2(new_n1139), .ZN(G381));
  NAND2_X1  g1036(.A1(new_n1188), .A2(new_n1214), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT122), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1188), .A2(new_n1187), .A3(new_n1214), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n673), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(new_n1238), .A2(new_n1239), .B1(new_n1240), .B2(new_n1185), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n1151), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1242), .A2(G384), .A3(G381), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n978), .A2(new_n1078), .A3(new_n1006), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1244), .A2(G396), .A3(G393), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1245), .ZN(G407));
  NAND2_X1  g1046(.A1(new_n644), .A2(G213), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(new_n1247), .B(KEYINPUT123), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(G407), .B(G213), .C1(new_n1242), .C2(new_n1249), .ZN(G409));
  XNOR2_X1  g1050(.A(new_n791), .B(G393), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT127), .ZN(new_n1252));
  AND3_X1   g1052(.A1(new_n978), .A2(new_n1006), .A3(new_n1078), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1078), .B1(new_n978), .B2(new_n1006), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1252), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G387), .A2(G390), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1256), .A2(KEYINPUT127), .A3(new_n1244), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1251), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1251), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1256), .A2(new_n1244), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1259), .B1(new_n1260), .B2(new_n1252), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1258), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT125), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT60), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(new_n1139), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT60), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(KEYINPUT125), .A3(new_n1149), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n673), .B1(new_n1269), .B2(KEYINPUT60), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1265), .A2(new_n1268), .A3(new_n1270), .ZN(new_n1271));
  AND3_X1   g1071(.A1(new_n1271), .A2(G384), .A3(new_n1234), .ZN(new_n1272));
  AOI21_X1  g1072(.A(G384), .B1(new_n1271), .B2(new_n1234), .ZN(new_n1273));
  OAI21_X1  g1073(.A(KEYINPUT126), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1271), .A2(new_n1234), .ZN(new_n1275));
  INV_X1    g1075(.A(G384), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT126), .ZN(new_n1278));
  NAND3_X1  g1078(.A1(new_n1271), .A2(G384), .A3(new_n1234), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1277), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1248), .A2(G2897), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1274), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1283), .A2(new_n1278), .A3(G2897), .A4(new_n1248), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1151), .B1(new_n1286), .B2(new_n1186), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1174), .A2(new_n1181), .A3(new_n1176), .A4(new_n940), .ZN(new_n1288));
  OAI21_X1  g1088(.A(KEYINPUT124), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT124), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1179), .A2(new_n1290), .A3(new_n1180), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1289), .A2(new_n730), .A3(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1151), .A2(new_n1288), .A3(new_n1214), .A4(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1249), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1285), .B1(new_n1287), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1294), .ZN(new_n1296));
  OAI211_X1 g1096(.A(new_n1296), .B(new_n1283), .C1(new_n1241), .C2(new_n1151), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT62), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(KEYINPUT62), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT61), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1262), .B1(new_n1298), .B2(new_n1301), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1300), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT63), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1303), .B1(new_n1304), .B2(new_n1297), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(G375), .A2(G378), .ZN(new_n1306));
  AOI22_X1  g1106(.A1(new_n1306), .A2(new_n1296), .B1(new_n1284), .B2(new_n1282), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1283), .ZN(new_n1308));
  AOI211_X1 g1108(.A(new_n1308), .B(new_n1294), .C1(G375), .C2(G378), .ZN(new_n1309));
  OAI21_X1  g1109(.A(KEYINPUT63), .B1(new_n1307), .B2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1305), .A2(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1302), .A2(new_n1311), .ZN(G405));
  NAND2_X1  g1112(.A1(new_n1242), .A2(new_n1306), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1283), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1242), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n1316), .B1(new_n1258), .B2(new_n1261), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1314), .A2(new_n1262), .A3(new_n1315), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1317), .A2(new_n1318), .ZN(G402));
endmodule


