//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n775, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  NOR2_X1   g000(.A1(G475), .A2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n192));
  NOR2_X1   g006(.A1(G125), .A2(G140), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(G125), .A2(G140), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n192), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G125), .ZN(new_n197));
  NOR3_X1   g011(.A1(new_n197), .A2(KEYINPUT16), .A3(G140), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n191), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n198), .ZN(new_n200));
  INV_X1    g014(.A(new_n195), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(new_n193), .ZN(new_n202));
  OAI211_X1 g016(.A(new_n200), .B(G146), .C1(new_n202), .C2(new_n192), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n199), .A2(KEYINPUT78), .A3(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT78), .ZN(new_n205));
  OAI211_X1 g019(.A(new_n205), .B(new_n191), .C1(new_n196), .C2(new_n198), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  NOR2_X1   g021(.A1(G237), .A2(G953), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G214), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT92), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n209), .A2(new_n210), .A3(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT92), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n212), .A2(new_n214), .A3(G214), .A4(new_n208), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n211), .A2(new_n215), .A3(KEYINPUT17), .A4(G131), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n211), .A2(new_n215), .ZN(new_n217));
  INV_X1    g031(.A(G131), .ZN(new_n218));
  XNOR2_X1  g032(.A(new_n217), .B(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n207), .B(new_n216), .C1(new_n219), .C2(KEYINPUT17), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT95), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT94), .B1(new_n211), .B2(new_n215), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT18), .A2(G131), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(new_n222), .B(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT93), .ZN(new_n226));
  INV_X1    g040(.A(new_n202), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n226), .B1(new_n227), .B2(new_n191), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT80), .B1(new_n194), .B2(new_n195), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT80), .ZN(new_n230));
  NOR3_X1   g044(.A1(new_n201), .A2(new_n193), .A3(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n191), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n202), .A2(KEYINPUT93), .A3(G146), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n228), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n221), .B1(new_n225), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT94), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n217), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n224), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n222), .A2(new_n223), .ZN(new_n239));
  AND4_X1   g053(.A1(new_n221), .A2(new_n234), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n190), .B(new_n220), .C1(new_n235), .C2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n234), .A2(new_n238), .A3(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT95), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n225), .A2(new_n221), .A3(new_n234), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n203), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT19), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n227), .A2(new_n248), .ZN(new_n249));
  OR2_X1    g063(.A1(new_n229), .A2(new_n231), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n250), .B2(new_n248), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n247), .B1(new_n251), .B2(new_n191), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n219), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n190), .B1(new_n246), .B2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n187), .B1(new_n242), .B2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT20), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT96), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n244), .A2(new_n245), .B1(new_n252), .B2(new_n219), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n241), .B(new_n258), .C1(new_n259), .C2(new_n190), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n253), .B1(new_n235), .B2(new_n240), .ZN(new_n262));
  INV_X1    g076(.A(new_n190), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n258), .B1(new_n264), .B2(new_n241), .ZN(new_n265));
  OAI211_X1 g079(.A(KEYINPUT20), .B(new_n187), .C1(new_n261), .C2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n246), .A2(new_n220), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n263), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n241), .ZN(new_n269));
  INV_X1    g083(.A(G902), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G475), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT99), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n213), .A2(G128), .ZN(new_n274));
  OR2_X1    g088(.A1(new_n274), .A2(KEYINPUT13), .ZN(new_n275));
  INV_X1    g089(.A(G128), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G143), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n277), .A3(KEYINPUT13), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n275), .A2(G134), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT97), .ZN(new_n280));
  INV_X1    g094(.A(G122), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G116), .ZN(new_n282));
  INV_X1    g096(.A(G116), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G122), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G107), .ZN(new_n286));
  INV_X1    g100(.A(G107), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n282), .A2(new_n284), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G134), .ZN(new_n289));
  XNOR2_X1  g103(.A(G128), .B(G143), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n286), .A2(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT97), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n275), .A2(new_n292), .A3(new_n278), .A4(G134), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n280), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT14), .B1(new_n281), .B2(G116), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT98), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT98), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n284), .A2(new_n297), .A3(KEYINPUT14), .ZN(new_n298));
  OR3_X1    g112(.A1(new_n281), .A2(KEYINPUT14), .A3(G116), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n296), .A2(new_n298), .A3(new_n299), .A4(new_n282), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G107), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n290), .B(new_n289), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n302), .A3(new_n288), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n273), .B1(new_n294), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  XOR2_X1   g119(.A(KEYINPUT9), .B(G234), .Z(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G217), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n307), .A2(new_n308), .A3(G953), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n294), .A2(new_n303), .A3(new_n273), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n305), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n309), .ZN(new_n312));
  INV_X1    g126(.A(new_n310), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n312), .B1(new_n313), .B2(new_n304), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n311), .A2(new_n314), .A3(new_n270), .ZN(new_n315));
  INV_X1    g129(.A(G478), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(KEYINPUT15), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(G234), .A2(G237), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(G902), .A3(G953), .ZN(new_n320));
  XOR2_X1   g134(.A(new_n320), .B(KEYINPUT100), .Z(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT21), .B(G898), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G953), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G952), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n325), .B1(G234), .B2(G237), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n323), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n317), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n311), .A2(new_n314), .A3(new_n270), .A4(new_n329), .ZN(new_n330));
  AND3_X1   g144(.A1(new_n318), .A2(new_n328), .A3(new_n330), .ZN(new_n331));
  AND4_X1   g145(.A1(new_n257), .A2(new_n266), .A3(new_n272), .A4(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(G214), .B1(G237), .B2(G902), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT2), .ZN(new_n335));
  INV_X1    g149(.A(G113), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(KEYINPUT68), .A2(KEYINPUT2), .A3(G113), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(KEYINPUT68), .B1(KEYINPUT2), .B2(G113), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n337), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(G116), .B(G119), .Z(new_n342));
  NOR3_X1   g156(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT70), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT70), .ZN(new_n344));
  NAND2_X1  g158(.A1(KEYINPUT2), .A2(G113), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT68), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  AOI22_X1  g161(.A1(new_n347), .A2(new_n338), .B1(new_n335), .B2(new_n336), .ZN(new_n348));
  XNOR2_X1  g162(.A(G116), .B(G119), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n344), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT69), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n342), .B1(new_n341), .B2(new_n351), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n348), .A2(KEYINPUT69), .ZN(new_n353));
  OAI22_X1  g167(.A1(new_n343), .A2(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT85), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n189), .A2(G107), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT3), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n189), .A2(G107), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT85), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n361), .B(KEYINPUT3), .C1(new_n189), .C2(G107), .ZN(new_n362));
  NAND4_X1  g176(.A1(new_n356), .A2(new_n359), .A3(new_n360), .A4(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G101), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n287), .A2(G104), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n358), .B2(new_n357), .ZN(new_n366));
  INV_X1    g180(.A(G101), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n366), .A2(new_n367), .A3(new_n356), .A4(new_n362), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n364), .A2(KEYINPUT4), .A3(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n363), .A2(new_n370), .A3(G101), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n354), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  OR3_X1    g186(.A1(new_n189), .A2(KEYINPUT86), .A3(G107), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n360), .A2(KEYINPUT86), .ZN(new_n374));
  OAI211_X1 g188(.A(new_n373), .B(G101), .C1(new_n374), .C2(new_n357), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n368), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT70), .B1(new_n341), .B2(new_n342), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n348), .A2(new_n344), .A3(new_n349), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n349), .A2(KEYINPUT5), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n283), .A2(KEYINPUT5), .A3(G119), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(new_n336), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n376), .A2(new_n379), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n372), .A2(new_n384), .ZN(new_n385));
  XOR2_X1   g199(.A(G110), .B(G122), .Z(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(new_n386), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n372), .A2(new_n384), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n387), .A2(KEYINPUT6), .A3(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n391), .A3(new_n386), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT65), .B1(new_n213), .B2(G146), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT65), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n191), .A3(G143), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT1), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n213), .A2(G146), .ZN(new_n398));
  NAND4_X1  g212(.A1(new_n396), .A2(new_n397), .A3(G128), .A4(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n213), .A2(G146), .ZN(new_n400));
  OAI21_X1  g214(.A(G128), .B1(new_n400), .B2(new_n397), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n191), .A2(G143), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(new_n398), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n399), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n197), .ZN(new_n406));
  OR2_X1    g220(.A1(KEYINPUT0), .A2(G128), .ZN(new_n407));
  NAND2_X1  g221(.A1(KEYINPUT0), .A2(G128), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n191), .A2(G143), .ZN(new_n409));
  OAI211_X1 g223(.A(new_n407), .B(new_n408), .C1(new_n400), .C2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT64), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n403), .A2(KEYINPUT64), .A3(new_n407), .A4(new_n408), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n396), .A2(KEYINPUT0), .A3(G128), .A4(new_n398), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n406), .B1(new_n197), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G224), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n417), .A2(G953), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n416), .B(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n390), .A2(new_n392), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT7), .B1(new_n417), .B2(G953), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n421), .A2(KEYINPUT91), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n416), .B(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n368), .A2(new_n375), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n379), .A2(new_n424), .A3(new_n383), .ZN(new_n425));
  XOR2_X1   g239(.A(new_n386), .B(KEYINPUT8), .Z(new_n426));
  XOR2_X1   g240(.A(new_n380), .B(KEYINPUT90), .Z(new_n427));
  AOI22_X1  g241(.A1(new_n427), .A2(new_n382), .B1(new_n378), .B2(new_n377), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n425), .B(new_n426), .C1(new_n428), .C2(new_n424), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n421), .A2(KEYINPUT91), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n423), .A2(new_n389), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n420), .A2(new_n431), .A3(new_n270), .ZN(new_n432));
  OAI21_X1  g246(.A(G210), .B1(G237), .B2(G902), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n420), .A2(new_n431), .A3(new_n270), .A4(new_n433), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n334), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XOR2_X1   g251(.A(KEYINPUT88), .B(G469), .Z(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n369), .A2(new_n415), .A3(new_n371), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT10), .ZN(new_n441));
  AOI211_X1 g255(.A(new_n276), .B(new_n409), .C1(new_n393), .C2(new_n395), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n396), .A2(new_n398), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n442), .A2(new_n397), .B1(new_n443), .B2(new_n401), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n441), .B1(new_n444), .B2(new_n424), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n399), .A2(new_n404), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n446), .A2(KEYINPUT10), .A3(new_n368), .A4(new_n375), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT11), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n289), .B2(G137), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n289), .A2(G137), .ZN(new_n450));
  INV_X1    g264(.A(G137), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(KEYINPUT11), .A3(G134), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G131), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n449), .A2(new_n452), .A3(new_n218), .A4(new_n450), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT87), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT87), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n454), .A2(new_n458), .A3(new_n455), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n440), .A2(new_n445), .A3(new_n447), .A4(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(G110), .B(G140), .ZN(new_n462));
  XNOR2_X1  g276(.A(new_n462), .B(KEYINPUT84), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n324), .A2(G227), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n463), .B(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n405), .A2(new_n424), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n444), .A2(new_n424), .ZN(new_n469));
  OAI211_X1 g283(.A(KEYINPUT12), .B(new_n456), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n456), .B1(new_n468), .B2(new_n469), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT12), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n466), .B1(new_n470), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n440), .A2(new_n445), .A3(new_n447), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(new_n456), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n465), .B1(new_n476), .B2(new_n461), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n270), .B(new_n439), .C1(new_n474), .C2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(G469), .A2(G902), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n461), .A2(new_n465), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n476), .ZN(new_n481));
  AND4_X1   g295(.A1(new_n440), .A2(new_n445), .A3(new_n447), .A4(new_n460), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n482), .B1(new_n473), .B2(new_n470), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n481), .B(G469), .C1(new_n483), .C2(new_n465), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n478), .A2(new_n479), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G221), .B1(new_n307), .B2(G902), .ZN(new_n486));
  AND3_X1   g300(.A1(new_n485), .A2(KEYINPUT89), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT89), .B1(new_n485), .B2(new_n486), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n332), .B(new_n437), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n451), .A2(G134), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n289), .A2(G137), .ZN(new_n492));
  OAI21_X1  g306(.A(G131), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n455), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT66), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n455), .A2(new_n493), .A3(KEYINPUT66), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n496), .A2(new_n446), .A3(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n456), .A2(new_n413), .A3(new_n412), .A4(new_n414), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT30), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(KEYINPUT67), .ZN(new_n503));
  INV_X1    g317(.A(new_n494), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n446), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(KEYINPUT30), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT67), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n500), .A2(new_n509), .A3(new_n501), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n503), .A2(new_n354), .A3(new_n508), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n341), .A2(new_n351), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n349), .B1(new_n348), .B2(KEYINPUT69), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n512), .A2(new_n513), .B1(new_n377), .B2(new_n378), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n499), .A3(new_n505), .ZN(new_n515));
  XOR2_X1   g329(.A(KEYINPUT26), .B(G101), .Z(new_n516));
  NAND2_X1  g330(.A1(new_n208), .A2(G210), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT72), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n515), .A2(new_n520), .A3(KEYINPUT72), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT31), .ZN(new_n526));
  AND3_X1   g340(.A1(new_n511), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n526), .B1(new_n511), .B2(new_n525), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT74), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n529), .B1(new_n499), .B2(new_n505), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n499), .A2(new_n529), .A3(new_n505), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n514), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT28), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XOR2_X1   g349(.A(KEYINPUT73), .B(KEYINPUT28), .Z(new_n536));
  INV_X1    g350(.A(new_n515), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n514), .B1(new_n499), .B2(new_n498), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n520), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  NOR3_X1   g354(.A1(new_n527), .A2(new_n528), .A3(new_n540), .ZN(new_n541));
  NOR2_X1   g355(.A1(G472), .A2(G902), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(KEYINPUT32), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n511), .A2(new_n525), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT31), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n535), .A2(new_n539), .ZN(new_n547));
  INV_X1    g361(.A(new_n520), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n511), .A2(new_n525), .A3(new_n526), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT32), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n551), .A2(new_n552), .A3(new_n542), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n507), .A2(new_n514), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT28), .B1(new_n554), .B2(new_n537), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n535), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n520), .A2(KEYINPUT29), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n270), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n511), .A2(new_n515), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n548), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT29), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n532), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n564), .A2(new_n530), .A3(new_n354), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n539), .B(new_n520), .C1(new_n565), .C2(KEYINPUT28), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT75), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT75), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n535), .A2(new_n568), .A3(new_n520), .A4(new_n539), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n559), .B1(new_n563), .B2(new_n570), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n544), .A2(new_n553), .B1(new_n571), .B2(G472), .ZN(new_n572));
  INV_X1    g386(.A(G234), .ZN(new_n573));
  OAI21_X1  g387(.A(G217), .B1(new_n573), .B2(G902), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(KEYINPUT76), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n324), .A2(G221), .A3(G234), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n576), .B(KEYINPUT22), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(G137), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n276), .A2(G119), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT77), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G119), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(G128), .ZN(new_n583));
  XOR2_X1   g397(.A(KEYINPUT24), .B(G110), .Z(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT23), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(G119), .B2(new_n276), .ZN(new_n587));
  NOR3_X1   g401(.A1(new_n582), .A2(KEYINPUT23), .A3(G128), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n583), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(G110), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n204), .A2(new_n206), .A3(new_n585), .A4(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(KEYINPUT79), .A2(G110), .ZN(new_n592));
  AND2_X1   g406(.A1(KEYINPUT79), .A2(G110), .ZN(new_n593));
  NOR3_X1   g407(.A1(new_n589), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n584), .B1(new_n581), .B2(new_n583), .ZN(new_n595));
  OAI211_X1 g409(.A(new_n232), .B(new_n203), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  AND3_X1   g410(.A1(new_n591), .A2(new_n596), .A3(KEYINPUT81), .ZN(new_n597));
  AOI21_X1  g411(.A(KEYINPUT81), .B1(new_n591), .B2(new_n596), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n578), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n578), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n591), .A2(new_n596), .ZN(new_n601));
  INV_X1    g415(.A(KEYINPUT81), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n599), .A2(new_n270), .A3(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT82), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT25), .ZN(new_n606));
  AND3_X1   g420(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n606), .B1(new_n604), .B2(new_n605), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n575), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n574), .A2(new_n270), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n599), .A2(new_n603), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NOR3_X1   g427(.A1(new_n572), .A2(KEYINPUT83), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT83), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n551), .A2(new_n552), .A3(new_n542), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n552), .B1(new_n551), .B2(new_n542), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n567), .A2(new_n569), .ZN(new_n618));
  AOI21_X1  g432(.A(KEYINPUT29), .B1(new_n560), .B2(new_n548), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n558), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(G472), .ZN(new_n621));
  OAI22_X1  g435(.A1(new_n616), .A2(new_n617), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n613), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n615), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n490), .B1(new_n614), .B2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(G101), .ZN(G3));
  NAND2_X1  g440(.A1(new_n551), .A2(new_n270), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n627), .A2(G472), .B1(new_n542), .B2(new_n551), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n628), .B(new_n623), .C1(new_n487), .C2(new_n488), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT101), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n485), .A2(new_n486), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT89), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n485), .A2(KEYINPUT89), .A3(new_n486), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n635), .A2(new_n636), .A3(new_n623), .A4(new_n628), .ZN(new_n637));
  AND2_X1   g451(.A1(new_n630), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n437), .A2(new_n328), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n266), .A2(new_n272), .A3(new_n257), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n311), .A2(new_n314), .A3(KEYINPUT102), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT33), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n311), .A2(new_n314), .A3(KEYINPUT102), .A4(KEYINPUT33), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(G478), .A3(new_n270), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n315), .A2(new_n316), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n640), .A2(new_n648), .ZN(new_n649));
  OAI21_X1  g463(.A(KEYINPUT103), .B1(new_n639), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n435), .A2(new_n436), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n651), .A2(new_n333), .A3(new_n328), .ZN(new_n652));
  INV_X1    g466(.A(new_n647), .ZN(new_n653));
  AOI21_X1  g467(.A(G902), .B1(new_n643), .B2(new_n644), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n653), .B1(new_n654), .B2(G478), .ZN(new_n655));
  INV_X1    g469(.A(new_n187), .ZN(new_n656));
  OAI21_X1  g470(.A(KEYINPUT96), .B1(new_n242), .B2(new_n254), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n656), .B1(new_n657), .B2(new_n260), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n658), .A2(KEYINPUT20), .B1(G475), .B2(new_n271), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n655), .B1(new_n659), .B2(new_n257), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT103), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n652), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n638), .A2(new_n650), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT34), .B(G104), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G6));
  OR2_X1    g479(.A1(new_n658), .A2(KEYINPUT20), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(new_n659), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n318), .A2(new_n330), .ZN(new_n668));
  INV_X1    g482(.A(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n639), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n638), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  NOR2_X1   g487(.A1(new_n600), .A2(KEYINPUT36), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT104), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n601), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n611), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n609), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n490), .A2(new_n628), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT105), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  INV_X1    g496(.A(G900), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n326), .B1(new_n321), .B2(new_n683), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n667), .A2(new_n669), .A3(new_n684), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n609), .A2(new_n677), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n544), .A2(new_n553), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n571), .A2(G472), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n686), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n651), .A2(new_n333), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n633), .B2(new_n634), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n685), .A2(new_n689), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G128), .ZN(G30));
  NAND2_X1  g507(.A1(new_n640), .A2(new_n668), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n684), .B(KEYINPUT39), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n695), .B1(new_n633), .B2(new_n634), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT40), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n694), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n651), .B(KEYINPUT38), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n554), .A2(new_n537), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n548), .A2(new_n702), .B1(new_n511), .B2(new_n525), .ZN(new_n703));
  OAI21_X1  g517(.A(G472), .B1(new_n703), .B2(G902), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n678), .B1(new_n687), .B2(new_n704), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n705), .B(new_n333), .C1(new_n696), .C2(new_n697), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n700), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(new_n213), .ZN(G45));
  INV_X1    g522(.A(new_n684), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n640), .A2(new_n648), .A3(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n689), .A2(new_n691), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT106), .B(G146), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G48));
  AOI21_X1  g527(.A(new_n613), .B1(new_n687), .B2(new_n688), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n270), .B1(new_n474), .B2(new_n477), .ZN(new_n715));
  OAI21_X1  g529(.A(G469), .B1(new_n715), .B2(KEYINPUT107), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n473), .A2(new_n470), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n480), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n476), .A2(new_n461), .ZN(new_n719));
  INV_X1    g533(.A(new_n465), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AOI21_X1  g535(.A(G902), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n486), .B(new_n478), .C1(new_n716), .C2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n662), .A2(new_n650), .A3(new_n714), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT41), .B(G113), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G15));
  NAND3_X1  g543(.A1(new_n670), .A2(new_n714), .A3(new_n726), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G116), .ZN(G18));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n725), .B2(new_n690), .ZN(new_n733));
  INV_X1    g547(.A(new_n478), .ZN(new_n734));
  INV_X1    g548(.A(G469), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n722), .B2(new_n723), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n715), .A2(KEYINPUT107), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n734), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(KEYINPUT108), .A3(new_n437), .A4(new_n486), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n332), .A3(new_n689), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(KEYINPUT109), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G119), .ZN(G21));
  AOI21_X1  g557(.A(new_n621), .B1(new_n551), .B2(new_n270), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n527), .A2(new_n528), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n556), .A2(new_n548), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n543), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n613), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n694), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n749), .A3(new_n652), .A4(new_n726), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G122), .ZN(G24));
  INV_X1    g565(.A(new_n744), .ZN(new_n752));
  INV_X1    g566(.A(new_n747), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n752), .A2(new_n678), .A3(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n640), .A2(new_n648), .A3(new_n709), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n740), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  XOR2_X1   g572(.A(new_n479), .B(KEYINPUT110), .Z(new_n759));
  AND3_X1   g573(.A1(new_n478), .A2(new_n484), .A3(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n486), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n334), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n651), .A2(new_n760), .A3(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n622), .A2(new_n710), .A3(new_n764), .A4(new_n623), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT42), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n714), .A2(KEYINPUT42), .A3(new_n710), .A4(new_n764), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT111), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT111), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n767), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G131), .ZN(G33));
  NAND3_X1  g588(.A1(new_n685), .A2(new_n714), .A3(new_n764), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G134), .ZN(G36));
  OAI21_X1  g590(.A(new_n481), .B1(new_n483), .B2(new_n465), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT45), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(G469), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n759), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT46), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(new_n478), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n761), .ZN(new_n783));
  INV_X1    g597(.A(new_n695), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT44), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n640), .A2(new_n655), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT43), .ZN(new_n787));
  INV_X1    g601(.A(new_n628), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n787), .A2(new_n788), .A3(new_n678), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n783), .B(new_n784), .C1(new_n785), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n785), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n435), .A2(new_n333), .A3(new_n436), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  OR2_X1    g608(.A1(new_n790), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G137), .ZN(G39));
  NAND2_X1  g610(.A1(new_n783), .A2(KEYINPUT47), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT47), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n782), .B2(new_n761), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n622), .A2(new_n623), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n800), .A2(new_n710), .A3(new_n793), .A4(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G140), .ZN(G42));
  NAND3_X1  g617(.A1(new_n786), .A2(new_n623), .A3(new_n762), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT112), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n687), .A2(new_n704), .ZN(new_n806));
  INV_X1    g620(.A(new_n699), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n738), .B(KEYINPUT49), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n805), .A2(new_n806), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n725), .A2(new_n327), .A3(new_n792), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n787), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n714), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(KEYINPUT48), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n787), .A2(new_n326), .A3(new_n748), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n738), .A2(new_n761), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n793), .B(new_n816), .C1(new_n800), .C2(new_n817), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n815), .A2(new_n333), .A3(new_n699), .A4(new_n725), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n819), .B(KEYINPUT50), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n806), .A2(new_n810), .A3(new_n623), .ZN(new_n821));
  OR3_X1    g635(.A1(new_n821), .A2(new_n640), .A3(new_n648), .ZN(new_n822));
  OR2_X1    g636(.A1(new_n811), .A2(new_n754), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n818), .A2(new_n820), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT51), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n814), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n813), .A2(KEYINPUT48), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n572), .A2(new_n667), .A3(new_n686), .A4(new_n668), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n792), .A2(new_n684), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n635), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(KEYINPUT113), .B1(new_n828), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n667), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n622), .A2(new_n833), .A3(new_n669), .A4(new_n678), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n834), .A2(new_n830), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n775), .B1(new_n832), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n649), .B1(new_n640), .B2(new_n669), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n630), .A2(new_n637), .A3(new_n652), .A4(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n756), .A2(new_n764), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n625), .A3(new_n679), .A4(new_n840), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n437), .B1(new_n487), .B2(new_n488), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n843), .A2(new_n572), .A3(new_n686), .ZN(new_n844));
  AOI22_X1  g658(.A1(new_n844), .A2(new_n685), .B1(new_n740), .B2(new_n756), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n437), .A2(new_n640), .A3(new_n668), .A4(new_n709), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n760), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n705), .A3(new_n486), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n845), .A2(KEYINPUT52), .A3(new_n711), .A4(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n757), .A2(new_n848), .A3(new_n692), .A4(new_n711), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n741), .A2(new_n727), .A3(new_n730), .A4(new_n750), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n854), .B1(new_n770), .B2(new_n772), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n842), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n856), .B(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT54), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n857), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT54), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n839), .A2(new_n625), .A3(new_n679), .ZN(new_n862));
  INV_X1    g676(.A(new_n775), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n828), .A2(KEYINPUT113), .A3(new_n831), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n835), .B1(new_n834), .B2(new_n830), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT114), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n862), .A2(new_n866), .A3(new_n867), .A4(new_n840), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT114), .B1(new_n837), .B2(new_n841), .ZN(new_n869));
  INV_X1    g683(.A(new_n769), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n870), .A2(new_n854), .A3(new_n857), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n868), .A2(new_n869), .A3(new_n853), .A4(new_n871), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n860), .A2(new_n861), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n826), .A2(new_n827), .A3(new_n859), .A4(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n824), .A2(new_n825), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n816), .A2(new_n740), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n325), .B(KEYINPUT115), .ZN(new_n878));
  OAI211_X1 g692(.A(new_n877), .B(new_n878), .C1(new_n649), .C2(new_n821), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n879), .B(KEYINPUT116), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n875), .A2(new_n876), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(G952), .A2(G953), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n809), .B1(new_n881), .B2(new_n882), .ZN(G75));
  AOI21_X1  g697(.A(new_n270), .B1(new_n860), .B2(new_n872), .ZN(new_n884));
  AOI21_X1  g698(.A(KEYINPUT56), .B1(new_n884), .B2(G210), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(KEYINPUT117), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n390), .A2(new_n392), .ZN(new_n887));
  XOR2_X1   g701(.A(new_n887), .B(new_n419), .Z(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT55), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n886), .B(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n324), .A2(G952), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n885), .A2(KEYINPUT117), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G51));
  INV_X1    g707(.A(KEYINPUT119), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n759), .B(KEYINPUT57), .Z(new_n895));
  AOI21_X1  g709(.A(new_n861), .B1(new_n860), .B2(new_n872), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n895), .B1(new_n873), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(KEYINPUT118), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT118), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n899), .B(new_n895), .C1(new_n873), .C2(new_n896), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n718), .A2(new_n721), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n894), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n902), .ZN(new_n904));
  AOI211_X1 g718(.A(KEYINPUT119), .B(new_n904), .C1(new_n898), .C2(new_n900), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n884), .A2(G469), .A3(new_n778), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n891), .B1(new_n906), .B2(new_n907), .ZN(G54));
  NAND3_X1  g722(.A1(new_n884), .A2(KEYINPUT58), .A3(G475), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n657), .A2(new_n260), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT120), .Z(new_n913));
  INV_X1    g727(.A(new_n891), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n909), .B2(new_n911), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n913), .A2(new_n915), .ZN(G60));
  XNOR2_X1  g730(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT122), .ZN(new_n918));
  NAND2_X1  g732(.A1(G478), .A2(G902), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n920), .B1(new_n643), .B2(new_n644), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n921), .B1(new_n873), .B2(new_n896), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n859), .B2(new_n874), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n914), .B(new_n922), .C1(new_n923), .C2(new_n645), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(G63));
  NAND2_X1  g739(.A1(new_n860), .A2(new_n872), .ZN(new_n926));
  NAND2_X1  g740(.A1(G217), .A2(G902), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n927), .B(KEYINPUT60), .Z(new_n928));
  NAND3_X1  g742(.A1(new_n926), .A2(new_n676), .A3(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT123), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n891), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n926), .A2(new_n928), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n599), .A2(new_n603), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT124), .ZN(new_n934));
  OAI221_X1 g748(.A(new_n931), .B1(new_n930), .B2(new_n929), .C1(new_n932), .C2(new_n934), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g750(.A(G953), .B1(new_n322), .B2(new_n417), .ZN(new_n937));
  INV_X1    g751(.A(new_n862), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(new_n854), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n939), .B2(G953), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n887), .B1(G898), .B2(new_n324), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n940), .B(new_n941), .ZN(G69));
  AOI21_X1  g756(.A(new_n324), .B1(G227), .B2(G900), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n812), .A2(new_n690), .A3(new_n694), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n783), .A2(new_n784), .A3(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n795), .A2(new_n711), .A3(new_n845), .A4(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n802), .A2(new_n773), .A3(new_n775), .ZN(new_n947));
  OR3_X1    g761(.A1(new_n946), .A2(new_n947), .A3(G953), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n503), .A2(new_n508), .A3(new_n510), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(new_n251), .Z(new_n950));
  OAI211_X1 g764(.A(new_n948), .B(new_n950), .C1(new_n683), .C2(new_n324), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n943), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n838), .A2(new_n793), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n954), .B(new_n696), .C1(new_n614), .C2(new_n624), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n955), .B1(new_n790), .B2(new_n794), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(KEYINPUT125), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT125), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n958), .B(new_n955), .C1(new_n790), .C2(new_n794), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n960), .A2(new_n802), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n845), .A2(new_n711), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n962), .A2(new_n707), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n963), .B(KEYINPUT62), .ZN(new_n964));
  AOI21_X1  g778(.A(G953), .B1(new_n961), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n951), .B1(new_n965), .B2(new_n950), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n953), .A2(new_n966), .ZN(new_n967));
  OAI221_X1 g781(.A(new_n951), .B1(new_n952), .B2(new_n943), .C1(new_n965), .C2(new_n950), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(G72));
  INV_X1    g783(.A(new_n560), .ZN(new_n970));
  NOR4_X1   g784(.A1(new_n946), .A2(new_n947), .A3(new_n938), .A4(new_n854), .ZN(new_n971));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT63), .Z(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n548), .B(new_n970), .C1(new_n971), .C2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n561), .A2(new_n545), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n858), .A2(new_n973), .A3(new_n976), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n977), .A2(new_n914), .ZN(new_n978));
  NAND4_X1  g792(.A1(new_n960), .A2(new_n802), .A3(new_n939), .A4(new_n964), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n973), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n980), .A2(new_n520), .A3(new_n560), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n975), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  INV_X1    g796(.A(KEYINPUT127), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(G57));
endmodule


