

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U553 ( .A(KEYINPUT29), .B(KEYINPUT94), .ZN(n701) );
  XNOR2_X1 U554 ( .A(n702), .B(n701), .ZN(n707) );
  NOR2_X1 U555 ( .A1(G164), .A2(G1384), .ZN(n792) );
  NOR2_X1 U556 ( .A1(G651), .A2(n637), .ZN(n648) );
  NOR2_X1 U557 ( .A1(G2104), .A2(G2105), .ZN(n519) );
  XOR2_X2 U558 ( .A(KEYINPUT17), .B(n519), .Z(n884) );
  NAND2_X1 U559 ( .A1(G138), .A2(n884), .ZN(n526) );
  INV_X1 U560 ( .A(G2105), .ZN(n520) );
  AND2_X1 U561 ( .A1(n520), .A2(G2104), .ZN(n883) );
  AND2_X1 U562 ( .A1(G102), .A2(n883), .ZN(n524) );
  NOR2_X1 U563 ( .A1(G2104), .A2(n520), .ZN(n887) );
  NAND2_X1 U564 ( .A1(G126), .A2(n887), .ZN(n522) );
  AND2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n888) );
  NAND2_X1 U566 ( .A1(G114), .A2(n888), .ZN(n521) );
  NAND2_X1 U567 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U568 ( .A1(n524), .A2(n523), .ZN(n525) );
  AND2_X1 U569 ( .A1(n526), .A2(n525), .ZN(G164) );
  NAND2_X1 U570 ( .A1(n884), .A2(G137), .ZN(n529) );
  NAND2_X1 U571 ( .A1(G101), .A2(n883), .ZN(n527) );
  XOR2_X1 U572 ( .A(n527), .B(KEYINPUT23), .Z(n528) );
  AND2_X1 U573 ( .A1(n529), .A2(n528), .ZN(n533) );
  NAND2_X1 U574 ( .A1(G125), .A2(n887), .ZN(n531) );
  NAND2_X1 U575 ( .A1(G113), .A2(n888), .ZN(n530) );
  AND2_X1 U576 ( .A1(n531), .A2(n530), .ZN(n532) );
  AND2_X1 U577 ( .A1(n533), .A2(n532), .ZN(G160) );
  AND2_X1 U578 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U579 ( .A(G57), .ZN(G237) );
  INV_X1 U580 ( .A(G82), .ZN(G220) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n637) );
  INV_X1 U582 ( .A(G651), .ZN(n537) );
  NOR2_X1 U583 ( .A1(n637), .A2(n537), .ZN(n640) );
  NAND2_X1 U584 ( .A1(G75), .A2(n640), .ZN(n536) );
  NOR2_X1 U585 ( .A1(G651), .A2(G543), .ZN(n534) );
  XOR2_X1 U586 ( .A(KEYINPUT65), .B(n534), .Z(n644) );
  NAND2_X1 U587 ( .A1(G88), .A2(n644), .ZN(n535) );
  NAND2_X1 U588 ( .A1(n536), .A2(n535), .ZN(n542) );
  NOR2_X1 U589 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X1 U590 ( .A(KEYINPUT1), .B(n538), .Z(n641) );
  NAND2_X1 U591 ( .A1(G62), .A2(n641), .ZN(n540) );
  NAND2_X1 U592 ( .A1(G50), .A2(n648), .ZN(n539) );
  NAND2_X1 U593 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U594 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U595 ( .A(KEYINPUT84), .B(n543), .Z(G303) );
  NAND2_X1 U596 ( .A1(G64), .A2(n641), .ZN(n545) );
  NAND2_X1 U597 ( .A1(G52), .A2(n648), .ZN(n544) );
  NAND2_X1 U598 ( .A1(n545), .A2(n544), .ZN(n551) );
  NAND2_X1 U599 ( .A1(n640), .A2(G77), .ZN(n546) );
  XOR2_X1 U600 ( .A(KEYINPUT67), .B(n546), .Z(n548) );
  NAND2_X1 U601 ( .A1(n644), .A2(G90), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U603 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U604 ( .A1(n551), .A2(n550), .ZN(G171) );
  NAND2_X1 U605 ( .A1(n644), .A2(G89), .ZN(n552) );
  XNOR2_X1 U606 ( .A(n552), .B(KEYINPUT4), .ZN(n554) );
  NAND2_X1 U607 ( .A1(G76), .A2(n640), .ZN(n553) );
  NAND2_X1 U608 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U609 ( .A(n555), .B(KEYINPUT5), .ZN(n561) );
  XNOR2_X1 U610 ( .A(KEYINPUT6), .B(KEYINPUT73), .ZN(n559) );
  NAND2_X1 U611 ( .A1(G63), .A2(n641), .ZN(n557) );
  NAND2_X1 U612 ( .A1(G51), .A2(n648), .ZN(n556) );
  NAND2_X1 U613 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U614 ( .A(n559), .B(n558), .ZN(n560) );
  NAND2_X1 U615 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U616 ( .A(KEYINPUT7), .B(n562), .ZN(G168) );
  XOR2_X1 U617 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U618 ( .A1(G7), .A2(G661), .ZN(n563) );
  XNOR2_X1 U619 ( .A(n563), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U620 ( .A(G223), .ZN(n824) );
  NAND2_X1 U621 ( .A1(n824), .A2(G567), .ZN(n564) );
  XOR2_X1 U622 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  XNOR2_X1 U623 ( .A(KEYINPUT13), .B(KEYINPUT71), .ZN(n570) );
  NAND2_X1 U624 ( .A1(G81), .A2(n644), .ZN(n565) );
  XNOR2_X1 U625 ( .A(n565), .B(KEYINPUT12), .ZN(n566) );
  XNOR2_X1 U626 ( .A(n566), .B(KEYINPUT70), .ZN(n568) );
  NAND2_X1 U627 ( .A1(G68), .A2(n640), .ZN(n567) );
  NAND2_X1 U628 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U629 ( .A(n570), .B(n569), .ZN(n573) );
  NAND2_X1 U630 ( .A1(n641), .A2(G56), .ZN(n571) );
  XOR2_X1 U631 ( .A(KEYINPUT14), .B(n571), .Z(n572) );
  NOR2_X1 U632 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U633 ( .A1(n648), .A2(G43), .ZN(n574) );
  NAND2_X1 U634 ( .A1(n575), .A2(n574), .ZN(n989) );
  INV_X1 U635 ( .A(G860), .ZN(n595) );
  OR2_X1 U636 ( .A1(n989), .A2(n595), .ZN(G153) );
  INV_X1 U637 ( .A(G171), .ZN(G301) );
  NAND2_X1 U638 ( .A1(G868), .A2(G301), .ZN(n585) );
  NAND2_X1 U639 ( .A1(G79), .A2(n640), .ZN(n577) );
  NAND2_X1 U640 ( .A1(G54), .A2(n648), .ZN(n576) );
  NAND2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n582) );
  NAND2_X1 U642 ( .A1(G92), .A2(n644), .ZN(n579) );
  NAND2_X1 U643 ( .A1(G66), .A2(n641), .ZN(n578) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(KEYINPUT72), .B(n580), .ZN(n581) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT15), .ZN(n975) );
  INV_X1 U648 ( .A(G868), .ZN(n651) );
  NAND2_X1 U649 ( .A1(n975), .A2(n651), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U651 ( .A1(G65), .A2(n641), .ZN(n587) );
  NAND2_X1 U652 ( .A1(G53), .A2(n648), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U654 ( .A(KEYINPUT68), .B(n588), .Z(n592) );
  NAND2_X1 U655 ( .A1(n640), .A2(G78), .ZN(n590) );
  NAND2_X1 U656 ( .A1(G91), .A2(n644), .ZN(n589) );
  AND2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U658 ( .A1(n592), .A2(n591), .ZN(G299) );
  NOR2_X1 U659 ( .A1(G286), .A2(n651), .ZN(n594) );
  NOR2_X1 U660 ( .A1(G868), .A2(G299), .ZN(n593) );
  NOR2_X1 U661 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U662 ( .A1(n595), .A2(G559), .ZN(n596) );
  INV_X1 U663 ( .A(n975), .ZN(n910) );
  NAND2_X1 U664 ( .A1(n596), .A2(n910), .ZN(n597) );
  XNOR2_X1 U665 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U666 ( .A1(G868), .A2(n989), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n910), .A2(G868), .ZN(n598) );
  NOR2_X1 U668 ( .A1(G559), .A2(n598), .ZN(n599) );
  NOR2_X1 U669 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U670 ( .A1(G123), .A2(n887), .ZN(n601) );
  XNOR2_X1 U671 ( .A(n601), .B(KEYINPUT74), .ZN(n602) );
  XNOR2_X1 U672 ( .A(KEYINPUT18), .B(n602), .ZN(n605) );
  NAND2_X1 U673 ( .A1(G135), .A2(n884), .ZN(n603) );
  XOR2_X1 U674 ( .A(KEYINPUT75), .B(n603), .Z(n604) );
  NAND2_X1 U675 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U676 ( .A1(G99), .A2(n883), .ZN(n607) );
  NAND2_X1 U677 ( .A1(G111), .A2(n888), .ZN(n606) );
  NAND2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n924) );
  XOR2_X1 U680 ( .A(G2096), .B(n924), .Z(n610) );
  NOR2_X1 U681 ( .A1(G2100), .A2(n610), .ZN(n611) );
  XOR2_X1 U682 ( .A(KEYINPUT76), .B(n611), .Z(G156) );
  NAND2_X1 U683 ( .A1(G55), .A2(n648), .ZN(n612) );
  XNOR2_X1 U684 ( .A(n612), .B(KEYINPUT78), .ZN(n619) );
  NAND2_X1 U685 ( .A1(G80), .A2(n640), .ZN(n614) );
  NAND2_X1 U686 ( .A1(G93), .A2(n644), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U688 ( .A1(G67), .A2(n641), .ZN(n615) );
  XNOR2_X1 U689 ( .A(KEYINPUT77), .B(n615), .ZN(n616) );
  NOR2_X1 U690 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n653) );
  NAND2_X1 U692 ( .A1(n910), .A2(G559), .ZN(n661) );
  XNOR2_X1 U693 ( .A(n989), .B(n661), .ZN(n620) );
  NOR2_X1 U694 ( .A1(G860), .A2(n620), .ZN(n621) );
  XOR2_X1 U695 ( .A(n653), .B(n621), .Z(G145) );
  NAND2_X1 U696 ( .A1(G73), .A2(n640), .ZN(n622) );
  XNOR2_X1 U697 ( .A(n622), .B(KEYINPUT2), .ZN(n630) );
  NAND2_X1 U698 ( .A1(G86), .A2(n644), .ZN(n624) );
  NAND2_X1 U699 ( .A1(G61), .A2(n641), .ZN(n623) );
  NAND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U701 ( .A(KEYINPUT82), .B(n625), .ZN(n628) );
  NAND2_X1 U702 ( .A1(G48), .A2(n648), .ZN(n626) );
  XNOR2_X1 U703 ( .A(KEYINPUT83), .B(n626), .ZN(n627) );
  NOR2_X1 U704 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(G305) );
  NAND2_X1 U706 ( .A1(n648), .A2(G49), .ZN(n631) );
  XNOR2_X1 U707 ( .A(KEYINPUT79), .B(n631), .ZN(n634) );
  NAND2_X1 U708 ( .A1(G651), .A2(G74), .ZN(n632) );
  XOR2_X1 U709 ( .A(KEYINPUT80), .B(n632), .Z(n633) );
  NOR2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n635) );
  XNOR2_X1 U711 ( .A(n635), .B(KEYINPUT81), .ZN(n636) );
  NOR2_X1 U712 ( .A1(n641), .A2(n636), .ZN(n639) );
  NAND2_X1 U713 ( .A1(n637), .A2(G87), .ZN(n638) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(G288) );
  NAND2_X1 U715 ( .A1(G72), .A2(n640), .ZN(n643) );
  NAND2_X1 U716 ( .A1(G60), .A2(n641), .ZN(n642) );
  NAND2_X1 U717 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U718 ( .A1(n644), .A2(G85), .ZN(n645) );
  XOR2_X1 U719 ( .A(KEYINPUT66), .B(n645), .Z(n646) );
  NOR2_X1 U720 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U721 ( .A1(n648), .A2(G47), .ZN(n649) );
  NAND2_X1 U722 ( .A1(n650), .A2(n649), .ZN(G290) );
  NAND2_X1 U723 ( .A1(n651), .A2(n653), .ZN(n652) );
  XNOR2_X1 U724 ( .A(n652), .B(KEYINPUT86), .ZN(n664) );
  XNOR2_X1 U725 ( .A(G303), .B(n653), .ZN(n660) );
  XNOR2_X1 U726 ( .A(G299), .B(G305), .ZN(n658) );
  XNOR2_X1 U727 ( .A(n989), .B(G288), .ZN(n656) );
  XNOR2_X1 U728 ( .A(KEYINPUT85), .B(KEYINPUT19), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n654), .B(G290), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n656), .B(n655), .ZN(n657) );
  XNOR2_X1 U731 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n660), .B(n659), .ZN(n909) );
  XNOR2_X1 U733 ( .A(n909), .B(n661), .ZN(n662) );
  NAND2_X1 U734 ( .A1(G868), .A2(n662), .ZN(n663) );
  NAND2_X1 U735 ( .A1(n664), .A2(n663), .ZN(G295) );
  NAND2_X1 U736 ( .A1(G2078), .A2(G2084), .ZN(n665) );
  XOR2_X1 U737 ( .A(KEYINPUT20), .B(n665), .Z(n666) );
  NAND2_X1 U738 ( .A1(G2090), .A2(n666), .ZN(n667) );
  XNOR2_X1 U739 ( .A(KEYINPUT21), .B(n667), .ZN(n668) );
  NAND2_X1 U740 ( .A1(n668), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U741 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U742 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U743 ( .A1(G220), .A2(G219), .ZN(n669) );
  XOR2_X1 U744 ( .A(KEYINPUT22), .B(n669), .Z(n670) );
  NOR2_X1 U745 ( .A1(G218), .A2(n670), .ZN(n671) );
  NAND2_X1 U746 ( .A1(G96), .A2(n671), .ZN(n831) );
  NAND2_X1 U747 ( .A1(n831), .A2(G2106), .ZN(n675) );
  NAND2_X1 U748 ( .A1(G69), .A2(G120), .ZN(n672) );
  NOR2_X1 U749 ( .A1(G237), .A2(n672), .ZN(n673) );
  NAND2_X1 U750 ( .A1(G108), .A2(n673), .ZN(n830) );
  NAND2_X1 U751 ( .A1(n830), .A2(G567), .ZN(n674) );
  NAND2_X1 U752 ( .A1(n675), .A2(n674), .ZN(n919) );
  NAND2_X1 U753 ( .A1(G483), .A2(G661), .ZN(n676) );
  NOR2_X1 U754 ( .A1(n919), .A2(n676), .ZN(n829) );
  NAND2_X1 U755 ( .A1(n829), .A2(G36), .ZN(G176) );
  AND2_X1 U756 ( .A1(G160), .A2(G40), .ZN(n677) );
  NAND2_X1 U757 ( .A1(n677), .A2(n792), .ZN(n678) );
  XNOR2_X2 U758 ( .A(KEYINPUT64), .B(n678), .ZN(n720) );
  INV_X1 U759 ( .A(n720), .ZN(n703) );
  NAND2_X1 U760 ( .A1(n703), .A2(G1996), .ZN(n679) );
  XNOR2_X1 U761 ( .A(n679), .B(KEYINPUT26), .ZN(n681) );
  NAND2_X1 U762 ( .A1(n720), .A2(G1341), .ZN(n680) );
  NAND2_X1 U763 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U764 ( .A1(n682), .A2(n989), .ZN(n686) );
  NAND2_X1 U765 ( .A1(G2067), .A2(n703), .ZN(n684) );
  NAND2_X1 U766 ( .A1(n720), .A2(G1348), .ZN(n683) );
  NAND2_X1 U767 ( .A1(n684), .A2(n683), .ZN(n687) );
  NOR2_X1 U768 ( .A1(n975), .A2(n687), .ZN(n685) );
  NOR2_X1 U769 ( .A1(n686), .A2(n685), .ZN(n689) );
  AND2_X1 U770 ( .A1(n975), .A2(n687), .ZN(n688) );
  NOR2_X1 U771 ( .A1(n689), .A2(n688), .ZN(n695) );
  INV_X1 U772 ( .A(G2072), .ZN(n950) );
  NOR2_X1 U773 ( .A1(n720), .A2(n950), .ZN(n691) );
  XNOR2_X1 U774 ( .A(KEYINPUT92), .B(KEYINPUT27), .ZN(n690) );
  XNOR2_X1 U775 ( .A(n691), .B(n690), .ZN(n693) );
  NAND2_X1 U776 ( .A1(n720), .A2(G1956), .ZN(n692) );
  NAND2_X1 U777 ( .A1(n693), .A2(n692), .ZN(n697) );
  NOR2_X1 U778 ( .A1(G299), .A2(n697), .ZN(n694) );
  NOR2_X1 U779 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U780 ( .A(KEYINPUT93), .B(n696), .ZN(n700) );
  NAND2_X1 U781 ( .A1(G299), .A2(n697), .ZN(n698) );
  XNOR2_X1 U782 ( .A(KEYINPUT28), .B(n698), .ZN(n699) );
  NAND2_X1 U783 ( .A1(n700), .A2(n699), .ZN(n702) );
  XOR2_X1 U784 ( .A(G2078), .B(KEYINPUT25), .Z(n951) );
  NAND2_X1 U785 ( .A1(n951), .A2(n703), .ZN(n705) );
  NAND2_X1 U786 ( .A1(n720), .A2(G1961), .ZN(n704) );
  NAND2_X1 U787 ( .A1(n705), .A2(n704), .ZN(n708) );
  NOR2_X1 U788 ( .A1(G301), .A2(n708), .ZN(n706) );
  NOR2_X1 U789 ( .A1(n707), .A2(n706), .ZN(n717) );
  NAND2_X1 U790 ( .A1(G301), .A2(n708), .ZN(n709) );
  XNOR2_X1 U791 ( .A(n709), .B(KEYINPUT95), .ZN(n714) );
  NAND2_X1 U792 ( .A1(n720), .A2(G8), .ZN(n766) );
  NOR2_X1 U793 ( .A1(G1966), .A2(n766), .ZN(n731) );
  NOR2_X1 U794 ( .A1(n720), .A2(G2084), .ZN(n732) );
  NOR2_X1 U795 ( .A1(n731), .A2(n732), .ZN(n710) );
  NAND2_X1 U796 ( .A1(G8), .A2(n710), .ZN(n711) );
  XNOR2_X1 U797 ( .A(KEYINPUT30), .B(n711), .ZN(n712) );
  NOR2_X1 U798 ( .A1(n712), .A2(G168), .ZN(n713) );
  NOR2_X1 U799 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U800 ( .A(n715), .B(KEYINPUT31), .ZN(n716) );
  NOR2_X1 U801 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U802 ( .A(n718), .B(KEYINPUT96), .ZN(n730) );
  INV_X1 U803 ( .A(n730), .ZN(n719) );
  AND2_X1 U804 ( .A1(n719), .A2(G286), .ZN(n728) );
  INV_X1 U805 ( .A(G8), .ZN(n726) );
  NOR2_X1 U806 ( .A1(n720), .A2(G2090), .ZN(n722) );
  NOR2_X1 U807 ( .A1(G1971), .A2(n766), .ZN(n721) );
  NOR2_X1 U808 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U809 ( .A1(G303), .A2(n723), .ZN(n724) );
  XOR2_X1 U810 ( .A(KEYINPUT97), .B(n724), .Z(n725) );
  NOR2_X1 U811 ( .A1(n726), .A2(n725), .ZN(n727) );
  NOR2_X1 U812 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U813 ( .A(n729), .B(KEYINPUT32), .ZN(n757) );
  NOR2_X1 U814 ( .A1(n731), .A2(n730), .ZN(n734) );
  NAND2_X1 U815 ( .A1(G8), .A2(n732), .ZN(n733) );
  NAND2_X1 U816 ( .A1(n734), .A2(n733), .ZN(n756) );
  NAND2_X1 U817 ( .A1(G288), .A2(G1976), .ZN(n735) );
  XOR2_X1 U818 ( .A(KEYINPUT98), .B(n735), .Z(n985) );
  NOR2_X1 U819 ( .A1(KEYINPUT99), .A2(n985), .ZN(n737) );
  INV_X1 U820 ( .A(n766), .ZN(n736) );
  NAND2_X1 U821 ( .A1(n737), .A2(n736), .ZN(n749) );
  INV_X1 U822 ( .A(n749), .ZN(n738) );
  AND2_X1 U823 ( .A1(n756), .A2(n738), .ZN(n745) );
  INV_X1 U824 ( .A(KEYINPUT99), .ZN(n740) );
  NOR2_X1 U825 ( .A1(G1976), .A2(G288), .ZN(n748) );
  NAND2_X1 U826 ( .A1(n748), .A2(KEYINPUT33), .ZN(n739) );
  NAND2_X1 U827 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U828 ( .A1(n748), .A2(KEYINPUT99), .ZN(n741) );
  NAND2_X1 U829 ( .A1(n742), .A2(n741), .ZN(n743) );
  NOR2_X1 U830 ( .A1(n766), .A2(n743), .ZN(n752) );
  INV_X1 U831 ( .A(n752), .ZN(n744) );
  AND2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U833 ( .A1(n757), .A2(n746), .ZN(n754) );
  NOR2_X1 U834 ( .A1(G303), .A2(G1971), .ZN(n747) );
  NOR2_X1 U835 ( .A1(n748), .A2(n747), .ZN(n987) );
  NOR2_X1 U836 ( .A1(n749), .A2(n987), .ZN(n750) );
  NOR2_X1 U837 ( .A1(n750), .A2(KEYINPUT33), .ZN(n751) );
  OR2_X1 U838 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U839 ( .A1(n754), .A2(n753), .ZN(n755) );
  XOR2_X1 U840 ( .A(G1981), .B(G305), .Z(n972) );
  NAND2_X1 U841 ( .A1(n755), .A2(n972), .ZN(n763) );
  NAND2_X1 U842 ( .A1(n757), .A2(n756), .ZN(n760) );
  NOR2_X1 U843 ( .A1(G2090), .A2(G303), .ZN(n758) );
  NAND2_X1 U844 ( .A1(G8), .A2(n758), .ZN(n759) );
  NAND2_X1 U845 ( .A1(n760), .A2(n759), .ZN(n761) );
  NAND2_X1 U846 ( .A1(n761), .A2(n766), .ZN(n762) );
  NAND2_X1 U847 ( .A1(n763), .A2(n762), .ZN(n812) );
  NOR2_X1 U848 ( .A1(G1981), .A2(G305), .ZN(n764) );
  XOR2_X1 U849 ( .A(n764), .B(KEYINPUT24), .Z(n765) );
  NOR2_X1 U850 ( .A1(n766), .A2(n765), .ZN(n810) );
  NAND2_X1 U851 ( .A1(n884), .A2(G141), .ZN(n767) );
  XNOR2_X1 U852 ( .A(KEYINPUT91), .B(n767), .ZN(n775) );
  NAND2_X1 U853 ( .A1(G129), .A2(n887), .ZN(n769) );
  NAND2_X1 U854 ( .A1(G117), .A2(n888), .ZN(n768) );
  NAND2_X1 U855 ( .A1(n769), .A2(n768), .ZN(n772) );
  NAND2_X1 U856 ( .A1(n883), .A2(G105), .ZN(n770) );
  XOR2_X1 U857 ( .A(KEYINPUT38), .B(n770), .Z(n771) );
  NOR2_X1 U858 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U859 ( .A(KEYINPUT90), .B(n773), .Z(n774) );
  OR2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n904) );
  NOR2_X1 U861 ( .A1(n904), .A2(G1996), .ZN(n776) );
  XNOR2_X1 U862 ( .A(n776), .B(KEYINPUT100), .ZN(n934) );
  INV_X1 U863 ( .A(G1991), .ZN(n947) );
  NAND2_X1 U864 ( .A1(n883), .A2(G95), .ZN(n779) );
  NAND2_X1 U865 ( .A1(G119), .A2(n887), .ZN(n777) );
  XOR2_X1 U866 ( .A(KEYINPUT89), .B(n777), .Z(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n783) );
  NAND2_X1 U868 ( .A1(G131), .A2(n884), .ZN(n781) );
  NAND2_X1 U869 ( .A1(G107), .A2(n888), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n782) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n895) );
  AND2_X1 U872 ( .A1(n947), .A2(n895), .ZN(n925) );
  NOR2_X1 U873 ( .A1(G1986), .A2(G290), .ZN(n784) );
  XOR2_X1 U874 ( .A(n784), .B(KEYINPUT101), .Z(n785) );
  NOR2_X1 U875 ( .A1(n925), .A2(n785), .ZN(n789) );
  NOR2_X1 U876 ( .A1(n895), .A2(n947), .ZN(n787) );
  AND2_X1 U877 ( .A1(n904), .A2(G1996), .ZN(n786) );
  NOR2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n920) );
  INV_X1 U879 ( .A(n920), .ZN(n788) );
  NOR2_X1 U880 ( .A1(n789), .A2(n788), .ZN(n790) );
  NOR2_X1 U881 ( .A1(n934), .A2(n790), .ZN(n791) );
  XNOR2_X1 U882 ( .A(n791), .B(KEYINPUT39), .ZN(n804) );
  NAND2_X1 U883 ( .A1(G160), .A2(G40), .ZN(n793) );
  NOR2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n814) );
  NAND2_X1 U885 ( .A1(G104), .A2(n883), .ZN(n795) );
  NAND2_X1 U886 ( .A1(G140), .A2(n884), .ZN(n794) );
  NAND2_X1 U887 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U888 ( .A(KEYINPUT34), .B(n796), .ZN(n801) );
  NAND2_X1 U889 ( .A1(G128), .A2(n887), .ZN(n798) );
  NAND2_X1 U890 ( .A1(G116), .A2(n888), .ZN(n797) );
  NAND2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n799) );
  XOR2_X1 U892 ( .A(n799), .B(KEYINPUT35), .Z(n800) );
  NOR2_X1 U893 ( .A1(n801), .A2(n800), .ZN(n802) );
  XOR2_X1 U894 ( .A(KEYINPUT36), .B(n802), .Z(n803) );
  XOR2_X1 U895 ( .A(KEYINPUT88), .B(n803), .Z(n903) );
  XNOR2_X1 U896 ( .A(G2067), .B(KEYINPUT37), .ZN(n805) );
  NOR2_X1 U897 ( .A1(n903), .A2(n805), .ZN(n923) );
  NAND2_X1 U898 ( .A1(n814), .A2(n923), .ZN(n816) );
  NAND2_X1 U899 ( .A1(n804), .A2(n816), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n903), .A2(n805), .ZN(n940) );
  NAND2_X1 U901 ( .A1(n806), .A2(n940), .ZN(n807) );
  XNOR2_X1 U902 ( .A(KEYINPUT102), .B(n807), .ZN(n808) );
  NAND2_X1 U903 ( .A1(n808), .A2(n814), .ZN(n820) );
  INV_X1 U904 ( .A(n820), .ZN(n809) );
  OR2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n811) );
  NOR2_X1 U906 ( .A1(n812), .A2(n811), .ZN(n822) );
  XNOR2_X1 U907 ( .A(KEYINPUT87), .B(G1986), .ZN(n813) );
  XNOR2_X1 U908 ( .A(n813), .B(G290), .ZN(n979) );
  NAND2_X1 U909 ( .A1(n979), .A2(n920), .ZN(n815) );
  AND2_X1 U910 ( .A1(n815), .A2(n814), .ZN(n818) );
  INV_X1 U911 ( .A(n816), .ZN(n817) );
  OR2_X1 U912 ( .A1(n818), .A2(n817), .ZN(n819) );
  AND2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n821) );
  NOR2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U915 ( .A(n823), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n824), .ZN(G217) );
  NAND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n826) );
  INV_X1 U918 ( .A(G661), .ZN(n825) );
  NOR2_X1 U919 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U920 ( .A(n827), .B(KEYINPUT105), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n828) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(G188) );
  INV_X1 U924 ( .A(G120), .ZN(G236) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G69), .ZN(G235) );
  NOR2_X1 U927 ( .A1(n831), .A2(n830), .ZN(n832) );
  XNOR2_X1 U928 ( .A(n832), .B(KEYINPUT106), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  XOR2_X1 U930 ( .A(G2454), .B(G2435), .Z(n834) );
  XNOR2_X1 U931 ( .A(G2438), .B(G2427), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n841) );
  XOR2_X1 U933 ( .A(KEYINPUT103), .B(G2446), .Z(n836) );
  XNOR2_X1 U934 ( .A(G2443), .B(G2430), .ZN(n835) );
  XNOR2_X1 U935 ( .A(n836), .B(n835), .ZN(n837) );
  XOR2_X1 U936 ( .A(n837), .B(G2451), .Z(n839) );
  XNOR2_X1 U937 ( .A(G1341), .B(G1348), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(n842) );
  NAND2_X1 U940 ( .A1(n842), .A2(G14), .ZN(n843) );
  XOR2_X1 U941 ( .A(KEYINPUT104), .B(n843), .Z(G401) );
  XOR2_X1 U942 ( .A(KEYINPUT109), .B(G1991), .Z(n845) );
  XNOR2_X1 U943 ( .A(G1996), .B(G1981), .ZN(n844) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U945 ( .A(n846), .B(G2474), .Z(n848) );
  XNOR2_X1 U946 ( .A(G1976), .B(G1986), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U948 ( .A(G1971), .B(G1956), .Z(n850) );
  XNOR2_X1 U949 ( .A(G1966), .B(G1961), .ZN(n849) );
  XNOR2_X1 U950 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U951 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U952 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n854), .B(n853), .ZN(G229) );
  XOR2_X1 U954 ( .A(KEYINPUT108), .B(KEYINPUT107), .Z(n856) );
  XNOR2_X1 U955 ( .A(G2678), .B(KEYINPUT43), .ZN(n855) );
  XNOR2_X1 U956 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U957 ( .A(KEYINPUT42), .B(G2090), .Z(n858) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2072), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U960 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U961 ( .A(G2096), .B(G2100), .ZN(n861) );
  XNOR2_X1 U962 ( .A(n862), .B(n861), .ZN(n864) );
  XOR2_X1 U963 ( .A(G2078), .B(G2084), .Z(n863) );
  XNOR2_X1 U964 ( .A(n864), .B(n863), .ZN(G227) );
  NAND2_X1 U965 ( .A1(n888), .A2(G112), .ZN(n865) );
  XOR2_X1 U966 ( .A(KEYINPUT111), .B(n865), .Z(n867) );
  NAND2_X1 U967 ( .A1(n883), .A2(G100), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U969 ( .A(KEYINPUT112), .B(n868), .ZN(n873) );
  NAND2_X1 U970 ( .A1(n887), .A2(G124), .ZN(n869) );
  XNOR2_X1 U971 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G136), .A2(n884), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U974 ( .A1(n873), .A2(n872), .ZN(G162) );
  NAND2_X1 U975 ( .A1(n883), .A2(G106), .ZN(n874) );
  XNOR2_X1 U976 ( .A(n874), .B(KEYINPUT114), .ZN(n876) );
  NAND2_X1 U977 ( .A1(G142), .A2(n884), .ZN(n875) );
  NAND2_X1 U978 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U979 ( .A(n877), .B(KEYINPUT45), .ZN(n882) );
  NAND2_X1 U980 ( .A1(G130), .A2(n887), .ZN(n879) );
  NAND2_X1 U981 ( .A1(G118), .A2(n888), .ZN(n878) );
  NAND2_X1 U982 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U983 ( .A(KEYINPUT113), .B(n880), .ZN(n881) );
  NAND2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n894) );
  NAND2_X1 U985 ( .A1(G103), .A2(n883), .ZN(n886) );
  NAND2_X1 U986 ( .A1(G139), .A2(n884), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n893) );
  NAND2_X1 U988 ( .A1(G127), .A2(n887), .ZN(n890) );
  NAND2_X1 U989 ( .A1(G115), .A2(n888), .ZN(n889) );
  NAND2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U991 ( .A(KEYINPUT47), .B(n891), .Z(n892) );
  NOR2_X1 U992 ( .A1(n893), .A2(n892), .ZN(n929) );
  XNOR2_X1 U993 ( .A(n894), .B(n929), .ZN(n899) );
  XOR2_X1 U994 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n897) );
  XNOR2_X1 U995 ( .A(G164), .B(n895), .ZN(n896) );
  XNOR2_X1 U996 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U997 ( .A(n899), .B(n898), .Z(n901) );
  XNOR2_X1 U998 ( .A(G160), .B(n924), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1000 ( .A(n902), .B(G162), .Z(n906) );
  XOR2_X1 U1001 ( .A(n904), .B(n903), .Z(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n907), .ZN(n908) );
  XOR2_X1 U1004 ( .A(KEYINPUT115), .B(n908), .Z(G395) );
  XOR2_X1 U1005 ( .A(n909), .B(G286), .Z(n912) );
  XNOR2_X1 U1006 ( .A(G171), .B(n910), .ZN(n911) );
  XNOR2_X1 U1007 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n913), .ZN(G397) );
  OR2_X1 U1009 ( .A1(n919), .A2(G401), .ZN(n916) );
  NOR2_X1 U1010 ( .A1(G229), .A2(G227), .ZN(n914) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n914), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(n916), .A2(n915), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n917) );
  NAND2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G303), .ZN(G166) );
  INV_X1 U1017 ( .A(n919), .ZN(G319) );
  INV_X1 U1018 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1019 ( .A(KEYINPUT117), .B(KEYINPUT52), .Z(n943) );
  XNOR2_X1 U1020 ( .A(G160), .B(G2084), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n927) );
  NOR2_X1 U1023 ( .A1(n925), .A2(n924), .ZN(n926) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(KEYINPUT116), .B(n928), .ZN(n939) );
  XOR2_X1 U1026 ( .A(G164), .B(G2078), .Z(n931) );
  XNOR2_X1 U1027 ( .A(n950), .B(n929), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(KEYINPUT50), .B(n932), .ZN(n937) );
  XOR2_X1 U1030 ( .A(G2090), .B(G162), .Z(n933) );
  NOR2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  XOR2_X1 U1032 ( .A(KEYINPUT51), .B(n935), .Z(n936) );
  NAND2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1036 ( .A(n943), .B(n942), .ZN(n944) );
  NOR2_X1 U1037 ( .A1(KEYINPUT55), .A2(n944), .ZN(n945) );
  XOR2_X1 U1038 ( .A(KEYINPUT118), .B(n945), .Z(n946) );
  NAND2_X1 U1039 ( .A1(n946), .A2(G29), .ZN(n1026) );
  XOR2_X1 U1040 ( .A(G29), .B(KEYINPUT122), .Z(n970) );
  XNOR2_X1 U1041 ( .A(G25), .B(n947), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n948), .A2(G28), .ZN(n949) );
  XNOR2_X1 U1043 ( .A(KEYINPUT119), .B(n949), .ZN(n961) );
  XNOR2_X1 U1044 ( .A(G33), .B(n950), .ZN(n955) );
  XNOR2_X1 U1045 ( .A(n951), .B(G27), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G1996), .B(G32), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n954) );
  NAND2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(KEYINPUT120), .B(G2067), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G26), .B(n956), .ZN(n957) );
  NOR2_X1 U1051 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1052 ( .A(KEYINPUT121), .B(n959), .Z(n960) );
  NAND2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(n962), .B(KEYINPUT53), .ZN(n965) );
  XOR2_X1 U1055 ( .A(G2084), .B(G34), .Z(n963) );
  XNOR2_X1 U1056 ( .A(KEYINPUT54), .B(n963), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n967) );
  XNOR2_X1 U1058 ( .A(G35), .B(G2090), .ZN(n966) );
  NOR2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(n968), .B(KEYINPUT55), .ZN(n969) );
  NAND2_X1 U1061 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n971), .ZN(n1024) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n995) );
  XNOR2_X1 U1064 ( .A(G1966), .B(G168), .ZN(n973) );
  NAND2_X1 U1065 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(n974), .B(KEYINPUT57), .ZN(n993) );
  XNOR2_X1 U1067 ( .A(G301), .B(G1961), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(n975), .B(G1348), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n983) );
  NAND2_X1 U1070 ( .A1(G303), .A2(G1971), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n979), .A2(n978), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G1956), .B(G299), .ZN(n980) );
  NOR2_X1 U1073 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1077 ( .A(KEYINPUT123), .B(n988), .Z(n991) );
  XNOR2_X1 U1078 ( .A(G1341), .B(n989), .ZN(n990) );
  NOR2_X1 U1079 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1080 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1081 ( .A1(n995), .A2(n994), .ZN(n1022) );
  INV_X1 U1082 ( .A(G16), .ZN(n1020) );
  XOR2_X1 U1083 ( .A(G1971), .B(G22), .Z(n998) );
  XOR2_X1 U1084 ( .A(G23), .B(KEYINPUT126), .Z(n996) );
  XNOR2_X1 U1085 ( .A(n996), .B(G1976), .ZN(n997) );
  NAND2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(G24), .B(G1986), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XOR2_X1 U1089 ( .A(KEYINPUT58), .B(n1001), .Z(n1017) );
  XOR2_X1 U1090 ( .A(G1961), .B(G5), .Z(n1012) );
  XOR2_X1 U1091 ( .A(G1348), .B(KEYINPUT59), .Z(n1002) );
  XNOR2_X1 U1092 ( .A(G4), .B(n1002), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G19), .B(G1341), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1008) );
  XNOR2_X1 U1095 ( .A(G1956), .B(G20), .ZN(n1006) );
  XNOR2_X1 U1096 ( .A(G6), .B(G1981), .ZN(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1098 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XOR2_X1 U1099 ( .A(KEYINPUT60), .B(n1009), .Z(n1010) );
  XNOR2_X1 U1100 ( .A(n1010), .B(KEYINPUT124), .ZN(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1102 ( .A(G21), .B(G1966), .ZN(n1013) );
  NOR2_X1 U1103 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1104 ( .A(KEYINPUT125), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(KEYINPUT61), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NAND2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NOR2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1110 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1111 ( .A(n1027), .B(KEYINPUT127), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(KEYINPUT62), .B(n1028), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

