

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785;

  BUF_X1 U368 ( .A(n657), .Z(n346) );
  NOR2_X1 U369 ( .A1(n445), .A2(G902), .ZN(n479) );
  INV_X2 U370 ( .A(G953), .ZN(n773) );
  NOR2_X2 U371 ( .A1(n353), .A2(n663), .ZN(n664) );
  NOR2_X2 U372 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U373 ( .A1(n448), .A2(n347), .ZN(n446) );
  NOR2_X2 U374 ( .A1(n611), .A2(KEYINPUT110), .ZN(n347) );
  XNOR2_X2 U375 ( .A(KEYINPUT91), .B(KEYINPUT90), .ZN(n554) );
  XNOR2_X2 U376 ( .A(G128), .B(G119), .ZN(n552) );
  AND2_X2 U377 ( .A1(n421), .A2(n364), .ZN(n420) );
  XOR2_X1 U378 ( .A(G116), .B(G119), .Z(n496) );
  XNOR2_X1 U379 ( .A(n477), .B(KEYINPUT39), .ZN(n634) );
  NOR2_X1 U380 ( .A1(n612), .A2(n611), .ZN(n348) );
  OR2_X1 U381 ( .A1(n387), .A2(KEYINPUT108), .ZN(n349) );
  NAND2_X2 U382 ( .A1(n656), .A2(n346), .ZN(n671) );
  AND2_X2 U383 ( .A1(n368), .A2(n694), .ZN(n371) );
  INV_X2 U384 ( .A(KEYINPUT23), .ZN(n372) );
  NOR2_X2 U385 ( .A1(n671), .A2(n659), .ZN(n661) );
  INV_X1 U386 ( .A(n657), .ZN(n586) );
  NAND2_X1 U387 ( .A1(n634), .A2(n360), .ZN(n467) );
  NOR2_X1 U388 ( .A1(n670), .A2(n611), .ZN(n587) );
  BUF_X1 U389 ( .A(n482), .Z(n354) );
  NOR2_X1 U390 ( .A1(n416), .A2(n355), .ZN(n415) );
  NAND2_X1 U391 ( .A1(n647), .A2(n651), .ZN(n611) );
  XNOR2_X1 U392 ( .A(n455), .B(G146), .ZN(n507) );
  INV_X1 U393 ( .A(G125), .ZN(n455) );
  NAND2_X1 U394 ( .A1(n370), .A2(n702), .ZN(n369) );
  NOR2_X1 U395 ( .A1(n637), .A2(n450), .ZN(n730) );
  AND2_X1 U396 ( .A1(n608), .A2(n607), .ZN(n382) );
  AND2_X1 U397 ( .A1(n386), .A2(n349), .ZN(n385) );
  NAND2_X1 U398 ( .A1(n415), .A2(n414), .ZN(n670) );
  XNOR2_X1 U399 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U400 ( .A(n488), .B(n499), .ZN(n487) );
  XNOR2_X1 U401 ( .A(n480), .B(n507), .ZN(n551) );
  INV_X1 U402 ( .A(n507), .ZN(n499) );
  XOR2_X1 U403 ( .A(G902), .B(KEYINPUT15), .Z(n695) );
  XOR2_X1 U404 ( .A(G113), .B(G104), .Z(n514) );
  XOR2_X1 U405 ( .A(G107), .B(G122), .Z(n524) );
  XNOR2_X1 U406 ( .A(KEYINPUT71), .B(G131), .ZN(n534) );
  NOR2_X1 U407 ( .A1(n351), .A2(n644), .ZN(n350) );
  XNOR2_X1 U408 ( .A(n624), .B(n483), .ZN(n351) );
  BUF_X1 U409 ( .A(n781), .Z(n352) );
  NOR2_X1 U410 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U411 ( .A(n624), .B(n483), .ZN(n645) );
  AND2_X2 U412 ( .A1(n463), .A2(n639), .ZN(n771) );
  XNOR2_X1 U413 ( .A(n350), .B(n485), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n646), .B(n485), .ZN(n679) );
  XNOR2_X1 U415 ( .A(n563), .B(n476), .ZN(n704) );
  XNOR2_X2 U416 ( .A(n454), .B(KEYINPUT22), .ZN(n656) );
  INV_X1 U417 ( .A(KEYINPUT0), .ZN(n485) );
  NOR2_X1 U418 ( .A1(G953), .A2(G237), .ZN(n538) );
  NAND2_X1 U419 ( .A1(n392), .A2(n389), .ZN(n388) );
  AND2_X1 U420 ( .A1(n360), .A2(n390), .ZN(n389) );
  OR2_X1 U421 ( .A1(n657), .A2(n393), .ZN(n392) );
  NOR2_X1 U422 ( .A1(G237), .A2(G902), .ZN(n505) );
  NAND2_X1 U423 ( .A1(n569), .A2(n437), .ZN(n436) );
  INV_X1 U424 ( .A(G902), .ZN(n437) );
  XNOR2_X1 U425 ( .A(n481), .B(KEYINPUT70), .ZN(n480) );
  INV_X1 U426 ( .A(KEYINPUT10), .ZN(n481) );
  XOR2_X1 U427 ( .A(G137), .B(G140), .Z(n565) );
  NAND2_X1 U428 ( .A1(n439), .A2(G902), .ZN(n438) );
  XNOR2_X1 U429 ( .A(n543), .B(n537), .ZN(n476) );
  XNOR2_X1 U430 ( .A(n541), .B(n452), .ZN(n543) );
  XNOR2_X1 U431 ( .A(n542), .B(n453), .ZN(n452) );
  AND2_X1 U432 ( .A1(n429), .A2(n484), .ZN(n425) );
  OR2_X1 U433 ( .A1(n357), .A2(n695), .ZN(n430) );
  NOR2_X1 U434 ( .A1(n419), .A2(n417), .ZN(n416) );
  XNOR2_X1 U435 ( .A(n513), .B(n410), .ZN(n744) );
  XNOR2_X1 U436 ( .A(n456), .B(n411), .ZN(n410) );
  INV_X1 U437 ( .A(G140), .ZN(n411) );
  XNOR2_X1 U438 ( .A(n769), .B(G146), .ZN(n535) );
  XNOR2_X1 U439 ( .A(G104), .B(G110), .ZN(n564) );
  XNOR2_X1 U440 ( .A(n376), .B(n375), .ZN(n463) );
  XNOR2_X1 U441 ( .A(n475), .B(KEYINPUT109), .ZN(n474) );
  INV_X1 U442 ( .A(n626), .ZN(n473) );
  INV_X1 U443 ( .A(KEYINPUT6), .ZN(n470) );
  AND2_X1 U444 ( .A1(n635), .A2(n444), .ZN(n625) );
  NAND2_X1 U445 ( .A1(n394), .A2(KEYINPUT107), .ZN(n393) );
  INV_X1 U446 ( .A(n623), .ZN(n394) );
  XNOR2_X1 U447 ( .A(G137), .B(G113), .ZN(n542) );
  INV_X1 U448 ( .A(KEYINPUT5), .ZN(n453) );
  XOR2_X1 U449 ( .A(KEYINPUT96), .B(KEYINPUT95), .Z(n540) );
  XNOR2_X1 U450 ( .A(n510), .B(n551), .ZN(n512) );
  XNOR2_X1 U451 ( .A(G122), .B(KEYINPUT98), .ZN(n508) );
  XOR2_X1 U452 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n509) );
  XNOR2_X1 U453 ( .A(n515), .B(n516), .ZN(n456) );
  XNOR2_X1 U454 ( .A(n534), .B(n533), .ZN(n769) );
  INV_X1 U455 ( .A(KEYINPUT72), .ZN(n532) );
  XNOR2_X1 U456 ( .A(n500), .B(n489), .ZN(n488) );
  XNOR2_X1 U457 ( .A(n504), .B(KEYINPUT17), .ZN(n489) );
  NAND2_X1 U458 ( .A1(n380), .A2(n377), .ZN(n376) );
  NOR2_X1 U459 ( .A1(n382), .A2(n381), .ZN(n380) );
  NAND2_X1 U460 ( .A1(n443), .A2(n441), .ZN(n381) );
  INV_X1 U461 ( .A(KEYINPUT48), .ZN(n375) );
  NAND2_X1 U462 ( .A1(G234), .A2(G237), .ZN(n491) );
  INV_X1 U463 ( .A(KEYINPUT38), .ZN(n449) );
  NAND2_X1 U464 ( .A1(n428), .A2(n359), .ZN(n427) );
  NAND2_X1 U465 ( .A1(n364), .A2(n423), .ZN(n422) );
  INV_X1 U466 ( .A(KEYINPUT28), .ZN(n413) );
  XNOR2_X1 U467 ( .A(n561), .B(n562), .ZN(n478) );
  XNOR2_X1 U468 ( .A(n372), .B(KEYINPUT89), .ZN(n555) );
  XNOR2_X1 U469 ( .A(G134), .B(G116), .ZN(n520) );
  NAND2_X1 U470 ( .A1(n384), .A2(n356), .ZN(n383) );
  INV_X1 U471 ( .A(KEYINPUT19), .ZN(n483) );
  XNOR2_X1 U472 ( .A(n517), .B(G475), .ZN(n518) );
  XNOR2_X1 U473 ( .A(n704), .B(n367), .ZN(n705) );
  XNOR2_X1 U474 ( .A(n744), .B(n366), .ZN(n745) );
  XNOR2_X1 U475 ( .A(n567), .B(n469), .ZN(n468) );
  INV_X1 U476 ( .A(G107), .ZN(n469) );
  XNOR2_X1 U477 ( .A(n566), .B(n490), .ZN(n567) );
  NOR2_X1 U478 ( .A1(G952), .A2(n773), .ZN(n756) );
  XNOR2_X1 U479 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U480 ( .A(n699), .B(KEYINPUT83), .ZN(n684) );
  XNOR2_X1 U481 ( .A(n472), .B(n471), .ZN(n637) );
  INV_X1 U482 ( .A(KEYINPUT43), .ZN(n471) );
  XNOR2_X1 U483 ( .A(n658), .B(KEYINPUT103), .ZN(n659) );
  INV_X1 U484 ( .A(KEYINPUT37), .ZN(n442) );
  AND2_X1 U485 ( .A1(n409), .A2(KEYINPUT1), .ZN(n355) );
  AND2_X1 U486 ( .A1(n387), .A2(KEYINPUT108), .ZN(n356) );
  INV_X1 U487 ( .A(KEYINPUT87), .ZN(n484) );
  AND2_X1 U488 ( .A1(n506), .A2(G210), .ZN(n357) );
  AND2_X1 U489 ( .A1(n432), .A2(n431), .ZN(n358) );
  OR2_X1 U490 ( .A1(n636), .A2(KEYINPUT87), .ZN(n359) );
  AND2_X1 U491 ( .A1(n617), .A2(n582), .ZN(n360) );
  AND2_X1 U492 ( .A1(n419), .A2(n417), .ZN(n361) );
  NAND2_X1 U493 ( .A1(n397), .A2(n398), .ZN(n362) );
  AND2_X1 U494 ( .A1(n771), .A2(KEYINPUT2), .ZN(n363) );
  INV_X1 U495 ( .A(n569), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n568), .B(G469), .ZN(n569) );
  AND2_X1 U497 ( .A1(n636), .A2(KEYINPUT87), .ZN(n364) );
  AND2_X1 U498 ( .A1(n771), .A2(n698), .ZN(n365) );
  INV_X1 U499 ( .A(KEYINPUT1), .ZN(n417) );
  INV_X1 U500 ( .A(KEYINPUT108), .ZN(n395) );
  XNOR2_X1 U501 ( .A(KEYINPUT59), .B(KEYINPUT67), .ZN(n366) );
  XNOR2_X1 U502 ( .A(KEYINPUT62), .B(KEYINPUT88), .ZN(n367) );
  NAND2_X1 U503 ( .A1(n697), .A2(n365), .ZN(n370) );
  XNOR2_X2 U504 ( .A(n403), .B(KEYINPUT45), .ZN(n697) );
  NAND2_X1 U505 ( .A1(n697), .A2(n363), .ZN(n368) );
  NAND2_X2 U506 ( .A1(n371), .A2(n369), .ZN(n703) );
  XNOR2_X1 U507 ( .A(n721), .B(n373), .ZN(n608) );
  INV_X1 U508 ( .A(KEYINPUT47), .ZN(n373) );
  XNOR2_X2 U509 ( .A(n374), .B(KEYINPUT81), .ZN(n721) );
  NAND2_X1 U510 ( .A1(n632), .A2(n640), .ZN(n374) );
  XNOR2_X1 U511 ( .A(n606), .B(KEYINPUT112), .ZN(n632) );
  XNOR2_X1 U512 ( .A(n379), .B(n378), .ZN(n377) );
  INV_X1 U513 ( .A(KEYINPUT46), .ZN(n378) );
  NAND2_X1 U514 ( .A1(n784), .A2(n785), .ZN(n379) );
  NAND2_X1 U515 ( .A1(n385), .A2(n383), .ZN(n635) );
  INV_X1 U516 ( .A(n388), .ZN(n384) );
  NAND2_X1 U517 ( .A1(n388), .A2(n395), .ZN(n386) );
  NAND2_X1 U518 ( .A1(n657), .A2(n391), .ZN(n387) );
  NAND2_X1 U519 ( .A1(n623), .A2(n391), .ZN(n390) );
  INV_X1 U520 ( .A(KEYINPUT107), .ZN(n391) );
  INV_X1 U521 ( .A(n675), .ZN(n396) );
  OR2_X2 U522 ( .A1(n740), .A2(n436), .ZN(n419) );
  INV_X1 U523 ( .A(n351), .ZN(n640) );
  NOR2_X1 U524 ( .A1(n672), .A2(n673), .ZN(n709) );
  NAND2_X1 U525 ( .A1(n651), .A2(n399), .ZN(n397) );
  OR2_X1 U526 ( .A1(n613), .A2(KEYINPUT110), .ZN(n398) );
  AND2_X1 U527 ( .A1(n647), .A2(n466), .ZN(n399) );
  NAND2_X1 U528 ( .A1(n418), .A2(n361), .ZN(n414) );
  NAND2_X1 U529 ( .A1(n435), .A2(n438), .ZN(n409) );
  BUF_X1 U530 ( .A(n780), .Z(n400) );
  BUF_X1 U531 ( .A(n663), .Z(n401) );
  XNOR2_X1 U532 ( .A(n433), .B(KEYINPUT35), .ZN(n780) );
  NAND2_X1 U533 ( .A1(n432), .A2(n431), .ZN(n421) );
  NOR2_X2 U534 ( .A1(n615), .A2(n616), .ZN(n629) );
  BUF_X1 U535 ( .A(n440), .Z(n402) );
  NAND2_X1 U536 ( .A1(n405), .A2(n404), .ZN(n403) );
  XNOR2_X1 U537 ( .A(n407), .B(KEYINPUT85), .ZN(n404) );
  NAND2_X1 U538 ( .A1(n406), .A2(n667), .ZN(n405) );
  XNOR2_X1 U539 ( .A(n666), .B(n662), .ZN(n406) );
  NAND2_X1 U540 ( .A1(n451), .A2(n683), .ZN(n407) );
  NOR2_X1 U541 ( .A1(n709), .A2(n682), .ZN(n683) );
  XNOR2_X1 U542 ( .A(n408), .B(n589), .ZN(n663) );
  NAND2_X1 U543 ( .A1(n586), .A2(n587), .ZN(n408) );
  NOR2_X2 U544 ( .A1(n465), .A2(n464), .ZN(n614) );
  INV_X1 U545 ( .A(n409), .ZN(n418) );
  OR2_X2 U546 ( .A1(n731), .A2(n430), .ZN(n429) );
  NAND2_X1 U547 ( .A1(n358), .A2(n425), .ZN(n424) );
  INV_X1 U548 ( .A(n612), .ZN(n448) );
  XOR2_X1 U549 ( .A(n622), .B(KEYINPUT82), .Z(n441) );
  XNOR2_X1 U550 ( .A(n519), .B(n518), .ZN(n582) );
  NOR2_X1 U551 ( .A1(n605), .A2(n412), .ZN(n606) );
  XNOR2_X1 U552 ( .A(n604), .B(n413), .ZN(n412) );
  NAND2_X2 U553 ( .A1(n418), .A2(n419), .ZN(n612) );
  NOR2_X1 U554 ( .A1(n420), .A2(n427), .ZN(n426) );
  OR2_X1 U555 ( .A1(n731), .A2(n422), .ZN(n428) );
  INV_X1 U556 ( .A(n430), .ZN(n423) );
  NAND2_X1 U557 ( .A1(n358), .A2(n429), .ZN(n450) );
  NAND2_X1 U558 ( .A1(n426), .A2(n424), .ZN(n624) );
  NAND2_X1 U559 ( .A1(n357), .A2(n695), .ZN(n431) );
  NAND2_X1 U560 ( .A1(n731), .A2(n357), .ZN(n432) );
  NAND2_X1 U561 ( .A1(n780), .A2(KEYINPUT44), .ZN(n668) );
  NAND2_X1 U562 ( .A1(n434), .A2(n665), .ZN(n433) );
  XNOR2_X1 U563 ( .A(n664), .B(KEYINPUT34), .ZN(n434) );
  NAND2_X1 U564 ( .A1(n740), .A2(n439), .ZN(n435) );
  OR2_X2 U565 ( .A1(n440), .A2(G101), .ZN(n502) );
  NAND2_X1 U566 ( .A1(n440), .A2(G101), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n402), .B(n770), .ZN(n775) );
  XNOR2_X2 U568 ( .A(n523), .B(KEYINPUT4), .ZN(n440) );
  XNOR2_X1 U569 ( .A(n443), .B(n442), .ZN(n727) );
  NAND2_X1 U570 ( .A1(n627), .A2(n626), .ZN(n443) );
  INV_X1 U571 ( .A(n624), .ZN(n444) );
  XNOR2_X1 U572 ( .A(n445), .B(n752), .ZN(n753) );
  XNOR2_X1 U573 ( .A(n559), .B(n768), .ZN(n445) );
  NAND2_X1 U574 ( .A1(n446), .A2(n362), .ZN(n465) );
  XNOR2_X1 U575 ( .A(n450), .B(n449), .ZN(n628) );
  AND2_X1 U576 ( .A1(n665), .A2(n450), .ZN(n620) );
  XNOR2_X1 U577 ( .A(n668), .B(KEYINPUT86), .ZN(n451) );
  NOR2_X2 U578 ( .A1(n679), .A2(n650), .ZN(n454) );
  XNOR2_X1 U579 ( .A(n459), .B(n457), .ZN(n558) );
  INV_X1 U580 ( .A(n458), .ZN(n457) );
  XNOR2_X1 U581 ( .A(n552), .B(n554), .ZN(n458) );
  XNOR2_X1 U582 ( .A(n553), .B(n555), .ZN(n459) );
  NAND2_X2 U583 ( .A1(n502), .A2(n503), .ZN(n536) );
  XNOR2_X1 U584 ( .A(n460), .B(n748), .ZN(G60) );
  NOR2_X2 U585 ( .A1(n747), .A2(n756), .ZN(n460) );
  XNOR2_X1 U586 ( .A(n461), .B(n708), .ZN(G57) );
  NOR2_X2 U587 ( .A1(n707), .A2(n756), .ZN(n461) );
  XNOR2_X1 U588 ( .A(n462), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U589 ( .A1(n736), .A2(n756), .ZN(n462) );
  AND2_X1 U590 ( .A1(n612), .A2(KEYINPUT110), .ZN(n464) );
  INV_X1 U591 ( .A(n613), .ZN(n466) );
  XNOR2_X2 U592 ( .A(n467), .B(n630), .ZN(n784) );
  XNOR2_X2 U593 ( .A(n563), .B(n468), .ZN(n740) );
  XNOR2_X2 U594 ( .A(n536), .B(n535), .ZN(n563) );
  XNOR2_X2 U595 ( .A(n677), .B(n470), .ZN(n657) );
  XNOR2_X2 U596 ( .A(n544), .B(n545), .ZN(n677) );
  NAND2_X1 U597 ( .A1(n474), .A2(n473), .ZN(n472) );
  NAND2_X1 U598 ( .A1(n635), .A2(n636), .ZN(n475) );
  NAND2_X1 U599 ( .A1(n629), .A2(n628), .ZN(n477) );
  XNOR2_X2 U600 ( .A(n479), .B(n478), .ZN(n651) );
  NAND2_X1 U601 ( .A1(n482), .A2(G472), .ZN(n706) );
  NAND2_X1 U602 ( .A1(n482), .A2(G210), .ZN(n735) );
  NAND2_X1 U603 ( .A1(n482), .A2(G475), .ZN(n746) );
  NAND2_X1 U604 ( .A1(n354), .A2(G469), .ZN(n741) );
  NAND2_X1 U605 ( .A1(n354), .A2(G478), .ZN(n749) );
  NAND2_X1 U606 ( .A1(n354), .A2(G217), .ZN(n754) );
  XNOR2_X2 U607 ( .A(n703), .B(KEYINPUT65), .ZN(n482) );
  XNOR2_X2 U608 ( .A(n486), .B(n762), .ZN(n731) );
  XNOR2_X2 U609 ( .A(n536), .B(n487), .ZN(n486) );
  XNOR2_X1 U610 ( .A(n498), .B(n497), .ZN(n762) );
  XNOR2_X2 U611 ( .A(n501), .B(G143), .ZN(n523) );
  XNOR2_X2 U612 ( .A(G128), .B(KEYINPUT64), .ZN(n501) );
  AND2_X1 U613 ( .A1(G227), .A2(n773), .ZN(n490) );
  XNOR2_X1 U614 ( .A(n532), .B(G134), .ZN(n533) );
  INV_X1 U615 ( .A(n537), .ZN(n497) );
  XNOR2_X1 U616 ( .A(n534), .B(KEYINPUT99), .ZN(n516) );
  INV_X1 U617 ( .A(n670), .ZN(n626) );
  INV_X1 U618 ( .A(n651), .ZN(n652) );
  INV_X1 U619 ( .A(KEYINPUT125), .ZN(n752) );
  NAND2_X1 U620 ( .A1(n473), .A2(n652), .ZN(n653) );
  XNOR2_X1 U621 ( .A(n706), .B(n705), .ZN(n707) );
  XNOR2_X1 U622 ( .A(n746), .B(n745), .ZN(n747) );
  XNOR2_X1 U623 ( .A(n754), .B(n753), .ZN(n755) );
  XNOR2_X1 U624 ( .A(n691), .B(n690), .ZN(G75) );
  XOR2_X1 U625 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n492) );
  XNOR2_X1 U626 ( .A(n492), .B(n491), .ZN(n600) );
  NAND2_X1 U627 ( .A1(G952), .A2(n600), .ZN(n599) );
  XOR2_X1 U628 ( .A(KEYINPUT16), .B(G110), .Z(n494) );
  XNOR2_X1 U629 ( .A(n524), .B(n514), .ZN(n493) );
  XNOR2_X1 U630 ( .A(n494), .B(n493), .ZN(n498) );
  XNOR2_X1 U631 ( .A(KEYINPUT3), .B(KEYINPUT74), .ZN(n495) );
  XNOR2_X1 U632 ( .A(n496), .B(n495), .ZN(n537) );
  NAND2_X1 U633 ( .A1(G224), .A2(n773), .ZN(n500) );
  INV_X1 U634 ( .A(KEYINPUT18), .ZN(n504) );
  XOR2_X1 U635 ( .A(KEYINPUT78), .B(n505), .Z(n506) );
  NAND2_X1 U636 ( .A1(n506), .A2(G214), .ZN(n636) );
  NAND2_X1 U637 ( .A1(n628), .A2(n636), .ZN(n583) );
  XNOR2_X1 U638 ( .A(n509), .B(n508), .ZN(n510) );
  NAND2_X1 U639 ( .A1(G214), .A2(n538), .ZN(n511) );
  XNOR2_X1 U640 ( .A(n512), .B(n511), .ZN(n513) );
  XNOR2_X1 U641 ( .A(G143), .B(n514), .ZN(n515) );
  NOR2_X1 U642 ( .A1(G902), .A2(n744), .ZN(n519) );
  XNOR2_X1 U643 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n517) );
  INV_X1 U644 ( .A(n582), .ZN(n618) );
  XOR2_X1 U645 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n521) );
  XNOR2_X1 U646 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U647 ( .A(n523), .B(n522), .ZN(n529) );
  XOR2_X1 U648 ( .A(n524), .B(KEYINPUT101), .Z(n527) );
  NAND2_X1 U649 ( .A1(G234), .A2(n773), .ZN(n525) );
  XOR2_X1 U650 ( .A(KEYINPUT8), .B(n525), .Z(n556) );
  NAND2_X1 U651 ( .A1(G217), .A2(n556), .ZN(n526) );
  XNOR2_X1 U652 ( .A(n527), .B(n526), .ZN(n528) );
  XNOR2_X1 U653 ( .A(n529), .B(n528), .ZN(n750) );
  NOR2_X1 U654 ( .A1(G902), .A2(n750), .ZN(n530) );
  XNOR2_X1 U655 ( .A(G478), .B(n530), .ZN(n617) );
  NAND2_X1 U656 ( .A1(n618), .A2(n617), .ZN(n649) );
  NOR2_X1 U657 ( .A1(n583), .A2(n649), .ZN(n531) );
  XOR2_X1 U658 ( .A(KEYINPUT41), .B(n531), .Z(n631) );
  INV_X1 U659 ( .A(n631), .ZN(n595) );
  XOR2_X1 U660 ( .A(KEYINPUT51), .B(KEYINPUT120), .Z(n579) );
  XNOR2_X1 U661 ( .A(G472), .B(KEYINPUT76), .ZN(n545) );
  NAND2_X1 U662 ( .A1(n538), .A2(G210), .ZN(n539) );
  XNOR2_X1 U663 ( .A(n540), .B(n539), .ZN(n541) );
  NOR2_X1 U664 ( .A1(n704), .A2(G902), .ZN(n544) );
  INV_X1 U665 ( .A(n677), .ZN(n609) );
  XOR2_X1 U666 ( .A(KEYINPUT94), .B(KEYINPUT21), .Z(n548) );
  INV_X1 U667 ( .A(n695), .ZN(n692) );
  NAND2_X1 U668 ( .A1(n692), .A2(G234), .ZN(n546) );
  XNOR2_X1 U669 ( .A(n546), .B(KEYINPUT20), .ZN(n560) );
  NAND2_X1 U670 ( .A1(n560), .A2(G221), .ZN(n547) );
  XNOR2_X1 U671 ( .A(n548), .B(n547), .ZN(n647) );
  XOR2_X1 U672 ( .A(KEYINPUT25), .B(KEYINPUT92), .Z(n550) );
  XNOR2_X1 U673 ( .A(KEYINPUT80), .B(KEYINPUT93), .ZN(n549) );
  XNOR2_X1 U674 ( .A(n550), .B(n549), .ZN(n562) );
  XNOR2_X1 U675 ( .A(n565), .B(n551), .ZN(n768) );
  XOR2_X1 U676 ( .A(KEYINPUT24), .B(G110), .Z(n553) );
  NAND2_X1 U677 ( .A1(G221), .A2(n556), .ZN(n557) );
  XNOR2_X1 U678 ( .A(n558), .B(n557), .ZN(n559) );
  NAND2_X1 U679 ( .A1(n560), .A2(G217), .ZN(n561) );
  XNOR2_X1 U680 ( .A(n565), .B(n564), .ZN(n566) );
  INV_X1 U681 ( .A(KEYINPUT73), .ZN(n568) );
  AND2_X1 U682 ( .A1(n609), .A2(n587), .ZN(n570) );
  XOR2_X1 U683 ( .A(KEYINPUT97), .B(n570), .Z(n674) );
  AND2_X1 U684 ( .A1(n611), .A2(n670), .ZN(n571) );
  XNOR2_X1 U685 ( .A(KEYINPUT50), .B(n571), .ZN(n576) );
  XNOR2_X1 U686 ( .A(KEYINPUT102), .B(n651), .ZN(n669) );
  NOR2_X1 U687 ( .A1(n647), .A2(n669), .ZN(n572) );
  XOR2_X1 U688 ( .A(KEYINPUT49), .B(n572), .Z(n573) );
  NOR2_X1 U689 ( .A1(n609), .A2(n573), .ZN(n574) );
  XNOR2_X1 U690 ( .A(KEYINPUT119), .B(n574), .ZN(n575) );
  NOR2_X1 U691 ( .A1(n576), .A2(n575), .ZN(n577) );
  NOR2_X1 U692 ( .A1(n674), .A2(n577), .ZN(n578) );
  XNOR2_X1 U693 ( .A(n579), .B(n578), .ZN(n580) );
  NOR2_X1 U694 ( .A1(n595), .A2(n580), .ZN(n592) );
  NOR2_X1 U695 ( .A1(n628), .A2(n636), .ZN(n581) );
  NOR2_X1 U696 ( .A1(n649), .A2(n581), .ZN(n585) );
  NOR2_X1 U697 ( .A1(n617), .A2(n582), .ZN(n724) );
  NOR2_X1 U698 ( .A1(n360), .A2(n724), .ZN(n681) );
  NOR2_X1 U699 ( .A1(n681), .A2(n583), .ZN(n584) );
  NOR2_X1 U700 ( .A1(n585), .A2(n584), .ZN(n590) );
  XOR2_X1 U701 ( .A(KEYINPUT33), .B(KEYINPUT75), .Z(n588) );
  XNOR2_X1 U702 ( .A(KEYINPUT105), .B(n588), .ZN(n589) );
  NOR2_X1 U703 ( .A1(n590), .A2(n401), .ZN(n591) );
  NOR2_X1 U704 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U705 ( .A(n593), .B(KEYINPUT52), .ZN(n594) );
  NOR2_X1 U706 ( .A1(n599), .A2(n594), .ZN(n598) );
  NOR2_X1 U707 ( .A1(n401), .A2(n595), .ZN(n596) );
  XOR2_X1 U708 ( .A(KEYINPUT121), .B(n596), .Z(n597) );
  NOR2_X1 U709 ( .A1(n598), .A2(n597), .ZN(n688) );
  NOR2_X1 U710 ( .A1(G953), .A2(n599), .ZN(n643) );
  NAND2_X1 U711 ( .A1(G902), .A2(n600), .ZN(n641) );
  OR2_X1 U712 ( .A1(n773), .A2(n641), .ZN(n601) );
  NOR2_X1 U713 ( .A1(G900), .A2(n601), .ZN(n602) );
  NOR2_X1 U714 ( .A1(n643), .A2(n602), .ZN(n613) );
  NOR2_X1 U715 ( .A1(n613), .A2(n651), .ZN(n603) );
  NAND2_X1 U716 ( .A1(n647), .A2(n603), .ZN(n623) );
  NOR2_X1 U717 ( .A1(n677), .A2(n623), .ZN(n604) );
  XOR2_X1 U718 ( .A(n612), .B(KEYINPUT111), .Z(n605) );
  NAND2_X1 U719 ( .A1(n721), .A2(n681), .ZN(n607) );
  NAND2_X1 U720 ( .A1(n681), .A2(KEYINPUT47), .ZN(n621) );
  NAND2_X1 U721 ( .A1(n636), .A2(n609), .ZN(n610) );
  XNOR2_X1 U722 ( .A(KEYINPUT30), .B(n610), .ZN(n616) );
  XNOR2_X1 U723 ( .A(n614), .B(KEYINPUT79), .ZN(n615) );
  OR2_X1 U724 ( .A1(n618), .A2(n617), .ZN(n619) );
  XOR2_X1 U725 ( .A(n619), .B(KEYINPUT106), .Z(n665) );
  NAND2_X1 U726 ( .A1(n629), .A2(n620), .ZN(n720) );
  NAND2_X1 U727 ( .A1(n621), .A2(n720), .ZN(n622) );
  XNOR2_X1 U728 ( .A(n625), .B(KEYINPUT36), .ZN(n627) );
  XOR2_X1 U729 ( .A(KEYINPUT113), .B(KEYINPUT40), .Z(n630) );
  NAND2_X1 U730 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U731 ( .A(n633), .B(KEYINPUT42), .ZN(n785) );
  NAND2_X1 U732 ( .A1(n724), .A2(n634), .ZN(n729) );
  INV_X1 U733 ( .A(n730), .ZN(n638) );
  AND2_X1 U734 ( .A1(n729), .A2(n638), .ZN(n639) );
  OR2_X1 U735 ( .A1(n773), .A2(G898), .ZN(n764) );
  NOR2_X1 U736 ( .A1(n641), .A2(n764), .ZN(n642) );
  NOR2_X1 U737 ( .A1(n643), .A2(n642), .ZN(n644) );
  INV_X1 U738 ( .A(n647), .ZN(n648) );
  OR2_X1 U739 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U740 ( .A1(n656), .A2(n677), .ZN(n654) );
  XNOR2_X1 U741 ( .A(n655), .B(KEYINPUT104), .ZN(n782) );
  NOR2_X1 U742 ( .A1(n473), .A2(n669), .ZN(n658) );
  XNOR2_X1 U743 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n660) );
  XNOR2_X1 U744 ( .A(n661), .B(n660), .ZN(n781) );
  NOR2_X2 U745 ( .A1(n782), .A2(n781), .ZN(n666) );
  INV_X1 U746 ( .A(KEYINPUT44), .ZN(n662) );
  NAND2_X1 U747 ( .A1(n666), .A2(n400), .ZN(n667) );
  NAND2_X1 U748 ( .A1(n670), .A2(n669), .ZN(n673) );
  XNOR2_X1 U749 ( .A(n671), .B(KEYINPUT84), .ZN(n672) );
  INV_X1 U750 ( .A(n353), .ZN(n675) );
  NAND2_X1 U751 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U752 ( .A(n676), .B(KEYINPUT31), .ZN(n725) );
  NAND2_X1 U753 ( .A1(n677), .A2(n348), .ZN(n678) );
  NOR2_X1 U754 ( .A1(n396), .A2(n678), .ZN(n711) );
  NOR2_X1 U755 ( .A1(n725), .A2(n711), .ZN(n680) );
  NOR2_X1 U756 ( .A1(n681), .A2(n680), .ZN(n682) );
  BUF_X1 U757 ( .A(n697), .Z(n757) );
  NAND2_X1 U758 ( .A1(n771), .A2(n757), .ZN(n685) );
  INV_X1 U759 ( .A(KEYINPUT2), .ZN(n699) );
  NOR2_X1 U760 ( .A1(G953), .A2(n686), .ZN(n687) );
  NAND2_X1 U761 ( .A1(n688), .A2(n687), .ZN(n691) );
  INV_X1 U762 ( .A(KEYINPUT122), .ZN(n689) );
  XNOR2_X1 U763 ( .A(n689), .B(KEYINPUT53), .ZN(n690) );
  INV_X1 U764 ( .A(KEYINPUT63), .ZN(n708) );
  OR2_X1 U765 ( .A1(KEYINPUT68), .A2(n692), .ZN(n693) );
  OR2_X1 U766 ( .A1(n699), .A2(n693), .ZN(n694) );
  INV_X1 U767 ( .A(KEYINPUT68), .ZN(n696) );
  OR2_X1 U768 ( .A1(n696), .A2(n695), .ZN(n698) );
  INV_X1 U769 ( .A(n698), .ZN(n701) );
  AND2_X1 U770 ( .A1(n699), .A2(KEYINPUT68), .ZN(n700) );
  OR2_X1 U771 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U772 ( .A(n709), .B(G101), .Z(G3) );
  NAND2_X1 U773 ( .A1(n711), .A2(n360), .ZN(n710) );
  XNOR2_X1 U774 ( .A(n710), .B(G104), .ZN(G6) );
  XNOR2_X1 U775 ( .A(G107), .B(KEYINPUT26), .ZN(n715) );
  XOR2_X1 U776 ( .A(KEYINPUT27), .B(KEYINPUT114), .Z(n713) );
  NAND2_X1 U777 ( .A1(n711), .A2(n724), .ZN(n712) );
  XNOR2_X1 U778 ( .A(n713), .B(n712), .ZN(n714) );
  XNOR2_X1 U779 ( .A(n715), .B(n714), .ZN(G9) );
  XOR2_X1 U780 ( .A(KEYINPUT29), .B(KEYINPUT117), .Z(n717) );
  NAND2_X1 U781 ( .A1(n721), .A2(n724), .ZN(n716) );
  XNOR2_X1 U782 ( .A(n717), .B(n716), .ZN(n719) );
  XOR2_X1 U783 ( .A(G128), .B(KEYINPUT116), .Z(n718) );
  XNOR2_X1 U784 ( .A(n719), .B(n718), .ZN(G30) );
  XNOR2_X1 U785 ( .A(G143), .B(n720), .ZN(G45) );
  NAND2_X1 U786 ( .A1(n721), .A2(n360), .ZN(n722) );
  XNOR2_X1 U787 ( .A(n722), .B(G146), .ZN(G48) );
  NAND2_X1 U788 ( .A1(n725), .A2(n360), .ZN(n723) );
  XNOR2_X1 U789 ( .A(n723), .B(G113), .ZN(G15) );
  NAND2_X1 U790 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U791 ( .A(n726), .B(G116), .ZN(G18) );
  XNOR2_X1 U792 ( .A(n727), .B(KEYINPUT118), .ZN(n728) );
  XNOR2_X1 U793 ( .A(G125), .B(n728), .ZN(G27) );
  XNOR2_X1 U794 ( .A(G134), .B(n729), .ZN(G36) );
  XOR2_X1 U795 ( .A(G140), .B(n730), .Z(G42) );
  BUF_X1 U796 ( .A(n731), .Z(n733) );
  XOR2_X1 U797 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n732) );
  XNOR2_X1 U798 ( .A(n735), .B(n734), .ZN(n736) );
  XOR2_X1 U799 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n738) );
  XNOR2_X1 U800 ( .A(KEYINPUT124), .B(KEYINPUT123), .ZN(n737) );
  XNOR2_X1 U801 ( .A(n738), .B(n737), .ZN(n739) );
  XOR2_X1 U802 ( .A(n740), .B(n739), .Z(n742) );
  XNOR2_X1 U803 ( .A(n742), .B(n741), .ZN(n743) );
  NOR2_X1 U804 ( .A1(n756), .A2(n743), .ZN(G54) );
  XOR2_X1 U805 ( .A(KEYINPUT60), .B(KEYINPUT69), .Z(n748) );
  XNOR2_X1 U806 ( .A(n750), .B(n749), .ZN(n751) );
  NOR2_X1 U807 ( .A1(n756), .A2(n751), .ZN(G63) );
  NOR2_X1 U808 ( .A1(n756), .A2(n755), .ZN(G66) );
  NAND2_X1 U809 ( .A1(n757), .A2(n773), .ZN(n761) );
  NAND2_X1 U810 ( .A1(G953), .A2(G224), .ZN(n758) );
  XNOR2_X1 U811 ( .A(KEYINPUT61), .B(n758), .ZN(n759) );
  NAND2_X1 U812 ( .A1(n759), .A2(G898), .ZN(n760) );
  NAND2_X1 U813 ( .A1(n761), .A2(n760), .ZN(n767) );
  XNOR2_X1 U814 ( .A(G101), .B(n762), .ZN(n763) );
  XNOR2_X1 U815 ( .A(n763), .B(KEYINPUT126), .ZN(n765) );
  NAND2_X1 U816 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U817 ( .A(n767), .B(n766), .Z(G69) );
  XNOR2_X1 U818 ( .A(n769), .B(n768), .ZN(n770) );
  XNOR2_X1 U819 ( .A(KEYINPUT127), .B(n775), .ZN(n772) );
  XNOR2_X1 U820 ( .A(n772), .B(n771), .ZN(n774) );
  NAND2_X1 U821 ( .A1(n774), .A2(n773), .ZN(n779) );
  XNOR2_X1 U822 ( .A(G227), .B(n775), .ZN(n776) );
  NAND2_X1 U823 ( .A1(n776), .A2(G900), .ZN(n777) );
  NAND2_X1 U824 ( .A1(n777), .A2(G953), .ZN(n778) );
  NAND2_X1 U825 ( .A1(n779), .A2(n778), .ZN(G72) );
  XOR2_X1 U826 ( .A(n400), .B(G122), .Z(G24) );
  XOR2_X1 U827 ( .A(n352), .B(G119), .Z(G21) );
  XNOR2_X1 U828 ( .A(G110), .B(KEYINPUT115), .ZN(n783) );
  XNOR2_X1 U829 ( .A(n783), .B(n782), .ZN(G12) );
  XNOR2_X1 U830 ( .A(n784), .B(G131), .ZN(G33) );
  XNOR2_X1 U831 ( .A(G137), .B(n785), .ZN(G39) );
endmodule

