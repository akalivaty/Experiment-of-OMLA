//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:37 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(G227gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT27), .B(G183gat), .ZN(new_n205));
  INV_X1    g004(.A(G190gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n208));
  XNOR2_X1  g007(.A(new_n207), .B(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(G169gat), .ZN(new_n210));
  INV_X1    g009(.A(G176gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT67), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT26), .ZN(new_n214));
  NOR2_X1   g013(.A1(G169gat), .A2(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT67), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n213), .A2(new_n214), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  AOI21_X1  g019(.A(new_n220), .B1(KEYINPUT26), .B2(new_n212), .ZN(new_n221));
  AOI22_X1  g020(.A1(new_n218), .A2(new_n221), .B1(G183gat), .B2(G190gat), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n209), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT23), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n212), .A2(new_n224), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n225), .A2(KEYINPUT25), .ZN(new_n226));
  XOR2_X1   g025(.A(new_n219), .B(KEYINPUT66), .Z(new_n227));
  INV_X1    g026(.A(KEYINPUT24), .ZN(new_n228));
  INV_X1    g027(.A(G183gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(new_n206), .ZN(new_n230));
  NAND3_X1  g029(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT68), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(new_n206), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT68), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n234), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n230), .A2(new_n232), .A3(new_n233), .A4(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n213), .A2(KEYINPUT23), .A3(new_n217), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n226), .A2(new_n227), .A3(new_n236), .A4(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n215), .A2(KEYINPUT23), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n225), .A2(new_n219), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT65), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(new_n229), .A3(new_n206), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT65), .B1(G183gat), .B2(G190gat), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n230), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT64), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n231), .B(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n240), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n238), .B1(new_n247), .B2(KEYINPUT25), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n238), .B(KEYINPUT69), .C1(new_n247), .C2(KEYINPUT25), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n223), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(KEYINPUT1), .ZN(new_n254));
  XNOR2_X1  g053(.A(G127gat), .B(G134gat), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT71), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259));
  INV_X1    g058(.A(G120gat), .ZN(new_n260));
  OR3_X1    g059(.A1(new_n257), .A2(new_n260), .A3(G113gat), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n258), .A2(new_n259), .A3(new_n255), .A4(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n252), .A2(new_n264), .ZN(new_n265));
  AOI211_X1 g064(.A(new_n263), .B(new_n223), .C1(new_n250), .C2(new_n251), .ZN(new_n266));
  OAI21_X1  g065(.A(new_n204), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT33), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT72), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n267), .A2(KEYINPUT72), .A3(new_n268), .ZN(new_n272));
  XNOR2_X1  g071(.A(G15gat), .B(G43gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(G71gat), .B(G99gat), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n275), .B1(new_n267), .B2(KEYINPUT32), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n271), .A2(new_n272), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT73), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT73), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n271), .A2(new_n279), .A3(new_n272), .A4(new_n276), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  OAI211_X1 g080(.A(new_n267), .B(KEYINPUT32), .C1(new_n268), .C2(new_n275), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  OR3_X1    g082(.A1(new_n265), .A2(new_n266), .A3(new_n204), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT34), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g085(.A(G78gat), .B(G106gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(G22gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT31), .B(G50gat), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT3), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n292));
  OR2_X1    g091(.A1(G197gat), .A2(G204gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(G197gat), .A2(G204gat), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n296));
  AND2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G211gat), .B(G218gat), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n295), .A2(new_n296), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n298), .B1(new_n297), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n291), .B1(new_n303), .B2(KEYINPUT29), .ZN(new_n304));
  XOR2_X1   g103(.A(G141gat), .B(G148gat), .Z(new_n305));
  XOR2_X1   g104(.A(G155gat), .B(G162gat), .Z(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(G155gat), .ZN(new_n308));
  INV_X1    g107(.A(G162gat), .ZN(new_n309));
  OAI21_X1  g108(.A(KEYINPUT2), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n305), .A2(new_n307), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n305), .A2(new_n310), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n306), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT77), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT77), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n304), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n311), .A2(new_n313), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n319), .B1(new_n320), .B2(KEYINPUT3), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n318), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n323), .A2(G228gat), .A3(G233gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n304), .A2(new_n320), .ZN(new_n325));
  NAND2_X1  g124(.A1(G228gat), .A2(G233gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n325), .A2(new_n326), .A3(new_n322), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n290), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n327), .A3(new_n290), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n288), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n330), .ZN(new_n332));
  INV_X1    g131(.A(new_n288), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n332), .A2(new_n333), .A3(new_n328), .ZN(new_n334));
  OR2_X1    g133(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n285), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n281), .A2(new_n337), .A3(new_n282), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n286), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n209), .A2(new_n222), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n248), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G226gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(new_n203), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n319), .B1(new_n343), .B2(new_n203), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n345), .B(new_n303), .C1(new_n252), .C2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G8gat), .B(G36gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G64gat), .B(G92gat), .ZN(new_n349));
  XOR2_X1   g148(.A(new_n348), .B(new_n349), .Z(new_n350));
  NOR2_X1   g149(.A1(new_n342), .A2(new_n346), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(new_n344), .B2(new_n252), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n347), .B(new_n350), .C1(new_n352), .C2(new_n303), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT30), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n347), .B1(new_n352), .B2(new_n303), .ZN(new_n357));
  INV_X1    g156(.A(new_n350), .ZN(new_n358));
  AOI22_X1  g157(.A1(new_n355), .A2(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n353), .A2(new_n356), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(KEYINPUT75), .ZN(new_n361));
  AND2_X1   g160(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G1gat), .B(G29gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT0), .ZN(new_n364));
  XNOR2_X1  g163(.A(G57gat), .B(G85gat), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n364), .B(new_n365), .Z(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n264), .A2(KEYINPUT4), .A3(new_n313), .A4(new_n311), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT4), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n263), .B2(new_n320), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G225gat), .A2(G233gat), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n291), .B1(new_n315), .B2(new_n316), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n263), .B1(new_n320), .B2(KEYINPUT3), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n372), .B(new_n373), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(new_n373), .ZN(new_n377));
  INV_X1    g176(.A(new_n316), .ZN(new_n378));
  OAI211_X1 g177(.A(KEYINPUT78), .B(new_n263), .C1(new_n378), .C2(new_n314), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n379), .B1(new_n263), .B2(new_n320), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n264), .B1(new_n315), .B2(new_n316), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(KEYINPUT78), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n377), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n376), .A2(new_n383), .A3(new_n384), .A4(KEYINPUT5), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n374), .A2(new_n375), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(new_n371), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT5), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n387), .A2(new_n388), .A3(new_n373), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n388), .B1(new_n387), .B2(new_n373), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n384), .B1(new_n391), .B2(new_n383), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n367), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n376), .A2(KEYINPUT5), .ZN(new_n394));
  INV_X1    g193(.A(new_n383), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT79), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n396), .A2(new_n366), .A3(new_n389), .A4(new_n385), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT6), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n393), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  OAI211_X1 g198(.A(KEYINPUT6), .B(new_n367), .C1(new_n390), .C2(new_n392), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  OR2_X1    g200(.A1(KEYINPUT83), .A2(KEYINPUT35), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n362), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n399), .A2(new_n400), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n359), .A2(new_n361), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n340), .B(new_n403), .C1(KEYINPUT83), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n339), .A2(KEYINPUT84), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n337), .B1(new_n281), .B2(new_n282), .ZN(new_n409));
  INV_X1    g208(.A(new_n282), .ZN(new_n410));
  AOI211_X1 g209(.A(new_n285), .B(new_n410), .C1(new_n278), .C2(new_n280), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n413), .A3(new_n336), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n403), .B1(new_n408), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT35), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n407), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AND2_X1   g216(.A1(new_n357), .A2(KEYINPUT37), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n358), .B1(new_n357), .B2(KEYINPUT37), .ZN(new_n419));
  OAI21_X1  g218(.A(KEYINPUT38), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n355), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n419), .A2(KEYINPUT38), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n352), .A2(new_n302), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n345), .B1(new_n252), .B2(new_n346), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT37), .B1(new_n425), .B2(new_n303), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT81), .ZN(new_n427));
  OR3_X1    g226(.A1(new_n424), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n427), .B1(new_n424), .B2(new_n426), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n421), .B1(new_n423), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT82), .B1(new_n404), .B2(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n428), .A2(new_n429), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n355), .B1(new_n433), .B2(new_n422), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT82), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n401), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n420), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n377), .B1(new_n386), .B2(new_n371), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n438), .A2(KEYINPUT80), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n438), .A2(KEYINPUT80), .ZN(new_n441));
  OR3_X1    g240(.A1(new_n380), .A2(new_n382), .A3(new_n377), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n440), .A2(KEYINPUT39), .A3(new_n441), .A4(new_n442), .ZN(new_n443));
  AND2_X1   g242(.A1(new_n440), .A2(new_n441), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n366), .B(new_n443), .C1(new_n444), .C2(KEYINPUT39), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT40), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n393), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n445), .A2(new_n446), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n335), .B1(new_n450), .B2(new_n405), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n437), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n412), .A2(KEYINPUT36), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT36), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n454), .B1(new_n409), .B2(new_n411), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n362), .A2(new_n401), .ZN(new_n456));
  AOI22_X1  g255(.A1(new_n453), .A2(new_n455), .B1(new_n335), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n417), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g258(.A(G15gat), .B(G22gat), .ZN(new_n460));
  OR2_X1    g259(.A1(new_n460), .A2(G1gat), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT88), .ZN(new_n462));
  AOI21_X1  g261(.A(G8gat), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT16), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n460), .B1(new_n464), .B2(G1gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g266(.A(new_n461), .B(new_n465), .C1(new_n462), .C2(G8gat), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(G50gat), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(G43gat), .ZN(new_n471));
  INV_X1    g270(.A(G43gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G50gat), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n471), .A2(new_n473), .A3(KEYINPUT15), .ZN(new_n474));
  NOR2_X1   g273(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n475));
  INV_X1    g274(.A(G36gat), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G29gat), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT86), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT86), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(G29gat), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n476), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g281(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n483));
  OAI211_X1 g282(.A(new_n474), .B(new_n477), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT17), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n471), .A2(new_n473), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT15), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n480), .A2(G29gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n478), .A2(KEYINPUT86), .ZN(new_n490));
  OAI21_X1  g289(.A(G36gat), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n471), .A2(new_n473), .A3(KEYINPUT15), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n488), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n483), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT87), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n477), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n475), .A2(KEYINPUT87), .A3(new_n476), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n484), .B(new_n485), .C1(new_n493), .C2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NOR4_X1   g299(.A1(new_n495), .A2(KEYINPUT14), .A3(G29gat), .A4(G36gat), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT87), .B1(new_n475), .B2(new_n476), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n483), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n503), .A2(new_n492), .A3(new_n488), .A4(new_n491), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n485), .B1(new_n504), .B2(new_n484), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n469), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(G229gat), .A2(G233gat), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n484), .B1(new_n493), .B2(new_n498), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n467), .A2(new_n468), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n506), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT18), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n506), .A2(KEYINPUT18), .A3(new_n507), .A4(new_n509), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n469), .A2(new_n504), .A3(new_n484), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n509), .ZN(new_n515));
  XOR2_X1   g314(.A(new_n507), .B(KEYINPUT13), .Z(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n512), .A2(new_n513), .A3(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT89), .ZN(new_n519));
  XNOR2_X1  g318(.A(G113gat), .B(G141gat), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(G197gat), .ZN(new_n521));
  XOR2_X1   g320(.A(KEYINPUT11), .B(G169gat), .Z(new_n522));
  XNOR2_X1  g321(.A(new_n521), .B(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT12), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n523), .A2(KEYINPUT12), .ZN(new_n526));
  NOR3_X1   g325(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT85), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT85), .ZN(new_n528));
  OR2_X1    g327(.A1(new_n523), .A2(KEYINPUT12), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n528), .B1(new_n529), .B2(new_n524), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n518), .A2(new_n519), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n524), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n512), .A2(new_n513), .A3(new_n517), .A4(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n519), .B1(new_n518), .B2(new_n531), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(G57gat), .A2(G64gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(G57gat), .A2(G64gat), .ZN(new_n541));
  OAI21_X1  g340(.A(KEYINPUT90), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(G57gat), .ZN(new_n543));
  INV_X1    g342(.A(G64gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT90), .ZN(new_n546));
  NAND2_X1  g345(.A1(G57gat), .A2(G64gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n542), .A2(new_n548), .A3(KEYINPUT9), .ZN(new_n549));
  AND2_X1   g348(.A1(G71gat), .A2(G78gat), .ZN(new_n550));
  NOR2_X1   g349(.A1(G71gat), .A2(G78gat), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT9), .ZN(new_n554));
  NOR3_X1   g353(.A1(new_n554), .A2(G71gat), .A3(G78gat), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n545), .B(new_n547), .C1(new_n555), .C2(new_n550), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n558), .A2(KEYINPUT21), .B1(new_n467), .B2(new_n468), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(KEYINPUT21), .ZN(new_n560));
  NAND2_X1  g359(.A1(G231gat), .A2(G233gat), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n560), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(G127gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n560), .B(new_n561), .ZN(new_n566));
  NOR2_X1   g365(.A1(new_n566), .A2(G127gat), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n559), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n566), .A2(G127gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n563), .A2(new_n564), .ZN(new_n570));
  INV_X1    g369(.A(new_n559), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(new_n308), .ZN(new_n575));
  XNOR2_X1  g374(.A(G183gat), .B(G211gat), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n575), .B(new_n576), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n568), .A2(new_n572), .A3(new_n577), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(G190gat), .B(G218gat), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n582), .B(KEYINPUT94), .Z(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(G99gat), .A2(G106gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT8), .ZN(new_n586));
  NAND2_X1  g385(.A1(G85gat), .A2(G92gat), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT7), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(G85gat), .ZN(new_n590));
  INV_X1    g389(.A(G92gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n593));
  NAND4_X1  g392(.A1(new_n586), .A2(new_n589), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G99gat), .B(G106gat), .ZN(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT92), .ZN(new_n598));
  AOI22_X1  g397(.A1(KEYINPUT8), .A2(new_n585), .B1(new_n590), .B2(new_n591), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n599), .A2(new_n595), .A3(new_n589), .A4(new_n593), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n597), .A2(new_n598), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n598), .B1(new_n597), .B2(new_n600), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g402(.A(KEYINPUT93), .B(new_n603), .C1(new_n500), .C2(new_n505), .ZN(new_n604));
  AND3_X1   g403(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n597), .A2(new_n600), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n605), .B1(new_n508), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n508), .A2(KEYINPUT17), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n499), .ZN(new_n611));
  AOI21_X1  g410(.A(KEYINPUT93), .B1(new_n611), .B2(new_n603), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n584), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT95), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G134gat), .B(G162gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT91), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n612), .ZN(new_n620));
  NAND4_X1  g419(.A1(new_n620), .A2(new_n583), .A3(new_n604), .A4(new_n608), .ZN(new_n621));
  AOI22_X1  g420(.A1(new_n615), .A2(new_n619), .B1(new_n613), .B2(new_n621), .ZN(new_n622));
  AND4_X1   g421(.A1(KEYINPUT95), .A2(new_n621), .A3(new_n613), .A4(new_n619), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n581), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(G120gat), .B(G148gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(G176gat), .B(G204gat), .ZN(new_n627));
  XOR2_X1   g426(.A(new_n626), .B(new_n627), .Z(new_n628));
  NAND2_X1  g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n553), .A2(new_n556), .B1(new_n600), .B2(new_n597), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n553), .A2(new_n600), .A3(new_n556), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT96), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n594), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n599), .A2(KEYINPUT96), .A3(new_n589), .A4(new_n593), .ZN(new_n635));
  AND3_X1   g434(.A1(new_n634), .A2(new_n596), .A3(new_n635), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n631), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n634), .A2(new_n596), .A3(new_n635), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n600), .A2(new_n556), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n638), .A2(new_n639), .A3(KEYINPUT97), .A4(new_n553), .ZN(new_n640));
  AOI211_X1 g439(.A(KEYINPUT10), .B(new_n630), .C1(new_n637), .C2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT10), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n557), .A2(new_n606), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n629), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n630), .ZN(new_n645));
  INV_X1    g444(.A(new_n552), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n545), .A2(new_n547), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n554), .B1(new_n647), .B2(KEYINPUT90), .ZN(new_n648));
  AOI21_X1  g447(.A(new_n646), .B1(new_n648), .B2(new_n548), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n600), .A2(new_n556), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(KEYINPUT97), .B1(new_n651), .B2(new_n638), .ZN(new_n652));
  AND4_X1   g451(.A1(KEYINPUT97), .A2(new_n638), .A3(new_n639), .A4(new_n553), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n645), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n629), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n628), .B1(new_n644), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n644), .A2(new_n656), .A3(new_n628), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n625), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT98), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT98), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n625), .A2(new_n664), .A3(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n459), .A2(new_n539), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g466(.A1(new_n667), .A2(new_n401), .ZN(new_n668));
  XOR2_X1   g467(.A(new_n668), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g468(.A1(new_n667), .A2(new_n362), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n670), .A2(KEYINPUT99), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(KEYINPUT99), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(G8gat), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT16), .B(G8gat), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n674), .B1(new_n671), .B2(new_n672), .ZN(new_n678));
  OAI211_X1 g477(.A(new_n673), .B(new_n677), .C1(new_n678), .C2(KEYINPUT42), .ZN(G1325gat));
  NAND2_X1  g478(.A1(new_n453), .A2(new_n455), .ZN(new_n680));
  OAI21_X1  g479(.A(G15gat), .B1(new_n667), .B2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n412), .ZN(new_n682));
  OR2_X1    g481(.A1(new_n682), .A2(G15gat), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n681), .B1(new_n667), .B2(new_n683), .ZN(G1326gat));
  NOR2_X1   g483(.A1(new_n667), .A2(new_n336), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT43), .B(G22gat), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  INV_X1    g486(.A(KEYINPUT45), .ZN(new_n688));
  INV_X1    g487(.A(new_n581), .ZN(new_n689));
  INV_X1    g488(.A(new_n539), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n689), .A2(new_n690), .A3(new_n660), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n459), .A2(new_n624), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n404), .A2(new_n479), .A3(new_n481), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n688), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  OR3_X1    g493(.A1(new_n692), .A2(new_n688), .A3(new_n693), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n403), .B1(new_n406), .B2(KEYINPUT83), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n696), .A2(new_n339), .ZN(new_n697));
  INV_X1    g496(.A(new_n403), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n413), .B1(new_n412), .B2(new_n336), .ZN(new_n699));
  NOR4_X1   g498(.A1(new_n409), .A2(new_n411), .A3(new_n335), .A4(KEYINPUT84), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n697), .B1(new_n701), .B2(KEYINPUT35), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n452), .A2(new_n457), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n624), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n459), .A2(KEYINPUT44), .A3(new_n624), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n706), .A2(new_n404), .A3(new_n707), .A4(new_n691), .ZN(new_n708));
  OAI22_X1  g507(.A1(new_n708), .A2(KEYINPUT100), .B1(new_n489), .B2(new_n490), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n708), .A2(KEYINPUT100), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n694), .B(new_n695), .C1(new_n709), .C2(new_n710), .ZN(G1328gat));
  NAND4_X1  g510(.A1(new_n706), .A2(new_n405), .A3(new_n707), .A4(new_n691), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n476), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n713), .B2(new_n712), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n692), .A2(G36gat), .A3(new_n362), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT46), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n715), .A2(new_n717), .ZN(G1329gat));
  AND2_X1   g517(.A1(new_n706), .A2(new_n707), .ZN(new_n719));
  INV_X1    g518(.A(new_n680), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n719), .A2(G43gat), .A3(new_n720), .A4(new_n691), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n459), .A2(new_n412), .A3(new_n624), .A4(new_n691), .ZN(new_n722));
  AOI22_X1  g521(.A1(new_n722), .A2(new_n472), .B1(KEYINPUT102), .B2(KEYINPUT47), .ZN(new_n723));
  OR2_X1    g522(.A1(KEYINPUT102), .A2(KEYINPUT47), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n721), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n721), .B2(new_n723), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(G1330gat));
  NAND4_X1  g526(.A1(new_n706), .A2(new_n335), .A3(new_n707), .A4(new_n691), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G50gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n335), .A2(new_n470), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n692), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n729), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT103), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT48), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n731), .B1(new_n728), .B2(G50gat), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT48), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n736), .A2(KEYINPUT103), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n735), .A2(new_n738), .ZN(G1331gat));
  NAND3_X1  g538(.A1(new_n625), .A2(new_n690), .A3(new_n660), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n740), .B(KEYINPUT104), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT105), .B1(new_n459), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n744));
  AOI211_X1 g543(.A(new_n744), .B(new_n741), .C1(new_n417), .C2(new_n458), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n404), .ZN(new_n747));
  XNOR2_X1  g546(.A(KEYINPUT106), .B(G57gat), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n747), .B(new_n748), .ZN(G1332gat));
  NOR2_X1   g548(.A1(new_n702), .A2(new_n703), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n744), .B1(new_n750), .B2(new_n741), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n459), .A2(KEYINPUT105), .A3(new_n742), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n362), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  AND2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n754), .B2(new_n755), .ZN(G1333gat));
  INV_X1    g557(.A(G71gat), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n753), .B2(new_n682), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n680), .A2(new_n759), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT107), .B1(new_n746), .B2(new_n761), .ZN(new_n762));
  AND4_X1   g561(.A1(KEYINPUT107), .A2(new_n751), .A3(new_n752), .A4(new_n761), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n760), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT50), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT50), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n766), .B(new_n760), .C1(new_n762), .C2(new_n763), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1334gat));
  NAND2_X1  g567(.A1(new_n746), .A2(new_n335), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g569(.A1(new_n689), .A2(new_n539), .A3(new_n661), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n706), .A2(new_n404), .A3(new_n707), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(G85gat), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n689), .A2(new_n539), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n459), .A2(new_n624), .A3(new_n774), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n661), .B1(new_n775), .B2(KEYINPUT51), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n776), .B1(KEYINPUT51), .B2(new_n775), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n404), .A2(new_n590), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n773), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(KEYINPUT108), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT108), .ZN(new_n781));
  OAI211_X1 g580(.A(new_n781), .B(new_n773), .C1(new_n777), .C2(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1336gat));
  NAND4_X1  g582(.A1(new_n706), .A2(new_n405), .A3(new_n707), .A4(new_n771), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G92gat), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n405), .A2(new_n591), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n777), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT52), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT52), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n789), .B(new_n785), .C1(new_n777), .C2(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(G1337gat));
  NAND3_X1  g590(.A1(new_n719), .A2(new_n720), .A3(new_n771), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(G99gat), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n682), .A2(G99gat), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n777), .B2(new_n794), .ZN(G1338gat));
  NAND4_X1  g594(.A1(new_n706), .A2(new_n335), .A3(new_n707), .A4(new_n771), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(G106gat), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n336), .A2(G106gat), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n797), .B1(new_n777), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT53), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT53), .ZN(new_n801));
  OAI211_X1 g600(.A(new_n801), .B(new_n797), .C1(new_n777), .C2(new_n798), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(G1339gat));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n643), .A2(new_n629), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT54), .B1(new_n641), .B2(new_n806), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n642), .B(new_n645), .C1(new_n652), .C2(new_n653), .ZN(new_n808));
  INV_X1    g607(.A(new_n643), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n655), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(KEYINPUT55), .B1(new_n807), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  OAI211_X1 g611(.A(new_n812), .B(new_n629), .C1(new_n641), .C2(new_n643), .ZN(new_n813));
  INV_X1    g612(.A(new_n628), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n804), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n628), .B1(new_n810), .B2(new_n812), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n812), .B1(new_n808), .B2(new_n805), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n644), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n817), .A2(new_n819), .A3(KEYINPUT109), .A4(KEYINPUT55), .ZN(new_n820));
  AND3_X1   g619(.A1(new_n816), .A2(new_n659), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n507), .B1(new_n506), .B2(new_n509), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT110), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n823), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n824), .B(new_n825), .C1(new_n515), .C2(new_n516), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(new_n523), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(new_n534), .ZN(new_n828));
  AOI21_X1  g627(.A(KEYINPUT55), .B1(new_n817), .B2(new_n819), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n829), .A2(new_n622), .A3(new_n623), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n821), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT111), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n660), .A2(new_n827), .A3(new_n534), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n819), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n535), .B2(new_n537), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n816), .A2(new_n659), .A3(new_n820), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n833), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n624), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT111), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n821), .A2(new_n828), .A3(new_n830), .A4(new_n842), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n832), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n581), .ZN(new_n845));
  NOR4_X1   g644(.A1(new_n581), .A2(new_n539), .A3(new_n624), .A4(new_n660), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT112), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n849));
  AOI211_X1 g648(.A(new_n849), .B(new_n846), .C1(new_n844), .C2(new_n581), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n851), .A2(new_n339), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n362), .A2(new_n404), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g654(.A(G113gat), .B1(new_n855), .B2(new_n690), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n856), .B(KEYINPUT113), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n851), .A2(new_n401), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n699), .A2(new_n700), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(new_n405), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n690), .A2(G113gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n857), .B1(new_n861), .B2(new_n862), .ZN(G1340gat));
  NOR3_X1   g662(.A1(new_n855), .A2(new_n260), .A3(new_n661), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n858), .A2(new_n660), .A3(new_n860), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n864), .B1(new_n260), .B2(new_n865), .ZN(G1341gat));
  OAI21_X1  g665(.A(G127gat), .B1(new_n855), .B2(new_n581), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n689), .A2(new_n564), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n867), .B1(new_n861), .B2(new_n868), .ZN(G1342gat));
  NOR3_X1   g668(.A1(new_n861), .A2(G134gat), .A3(new_n840), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  OR2_X1    g670(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n872));
  OAI21_X1  g671(.A(G134gat), .B1(new_n855), .B2(new_n840), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(KEYINPUT56), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G1343gat));
  NAND2_X1  g674(.A1(new_n680), .A2(new_n335), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n876), .A2(new_n405), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n858), .A2(new_n877), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n878), .A2(G141gat), .A3(new_n690), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n879), .A2(KEYINPUT58), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n881));
  AOI22_X1  g680(.A1(KEYINPUT111), .A2(new_n831), .B1(new_n839), .B2(new_n840), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n689), .B1(new_n882), .B2(new_n843), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n849), .B1(new_n883), .B2(new_n846), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n845), .A2(KEYINPUT112), .A3(new_n847), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n336), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n881), .B1(new_n886), .B2(KEYINPUT57), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n335), .B1(new_n848), .B2(new_n850), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n888), .A2(KEYINPUT114), .A3(new_n889), .ZN(new_n890));
  AOI211_X1 g689(.A(new_n889), .B(new_n336), .C1(new_n845), .C2(new_n847), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n887), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n680), .A2(new_n854), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n893), .A2(new_n539), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT116), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G141gat), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n896), .A2(KEYINPUT116), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n880), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n896), .A2(KEYINPUT115), .A3(G141gat), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT115), .B1(new_n896), .B2(G141gat), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n901), .A2(new_n902), .A3(new_n879), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(G1344gat));
  INV_X1    g704(.A(G148gat), .ZN(new_n906));
  AND4_X1   g705(.A1(new_n906), .A2(new_n858), .A3(new_n660), .A4(new_n877), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT117), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n666), .A2(new_n690), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n821), .A2(new_n830), .A3(KEYINPUT119), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n828), .ZN(new_n911));
  AOI21_X1  g710(.A(KEYINPUT119), .B1(new_n821), .B2(new_n830), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n841), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(new_n581), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n909), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n336), .A2(KEYINPUT57), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n888), .A2(KEYINPUT57), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n894), .A2(new_n661), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n906), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT120), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n915), .A2(new_n916), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n922), .B1(new_n886), .B2(new_n889), .ZN(new_n923));
  INV_X1    g722(.A(new_n918), .ZN(new_n924));
  OAI21_X1  g723(.A(G148gat), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n926));
  INV_X1    g725(.A(new_n920), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n925), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n921), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g728(.A1(new_n906), .A2(KEYINPUT59), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n888), .A2(new_n889), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n891), .B1(new_n931), .B2(new_n881), .ZN(new_n932));
  AOI21_X1  g731(.A(new_n894), .B1(new_n932), .B2(new_n890), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n930), .B1(new_n933), .B2(new_n660), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n908), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT121), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n908), .B(new_n937), .C1(new_n929), .C2(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1345gat));
  INV_X1    g738(.A(new_n878), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n940), .A2(new_n308), .A3(new_n689), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n933), .A2(new_n689), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n941), .B1(new_n942), .B2(new_n308), .ZN(G1346gat));
  AOI21_X1  g742(.A(G162gat), .B1(new_n940), .B2(new_n624), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n840), .A2(new_n309), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n944), .B1(new_n933), .B2(new_n945), .ZN(G1347gat));
  NOR2_X1   g745(.A1(new_n362), .A2(new_n404), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NOR3_X1   g747(.A1(new_n851), .A2(new_n339), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n210), .B1(new_n949), .B2(new_n539), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT123), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n401), .B1(new_n848), .B2(new_n850), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n953));
  XNOR2_X1  g752(.A(new_n952), .B(new_n953), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n859), .A2(new_n362), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n539), .A2(new_n210), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(G1348gat));
  INV_X1    g757(.A(new_n949), .ZN(new_n959));
  OAI21_X1  g758(.A(G176gat), .B1(new_n959), .B2(new_n661), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n660), .A2(new_n211), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n960), .B1(new_n956), .B2(new_n961), .ZN(G1349gat));
  NAND2_X1  g761(.A1(new_n689), .A2(new_n205), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n959), .A2(new_n581), .ZN(new_n964));
  OAI22_X1  g763(.A1(new_n956), .A2(new_n963), .B1(new_n229), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT60), .ZN(G1350gat));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n624), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(new_n968), .A3(G190gat), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n968), .B1(new_n967), .B2(G190gat), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n624), .A2(new_n206), .ZN(new_n972));
  OAI22_X1  g771(.A1(new_n970), .A2(new_n971), .B1(new_n956), .B2(new_n972), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT124), .ZN(G1351gat));
  NOR3_X1   g773(.A1(new_n923), .A2(new_n720), .A3(new_n948), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(G197gat), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n976), .A2(new_n977), .A3(new_n690), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n876), .A2(new_n362), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n954), .A2(new_n979), .ZN(new_n980));
  OR2_X1    g779(.A1(new_n980), .A2(KEYINPUT125), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(KEYINPUT125), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n981), .A2(new_n539), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n978), .B1(new_n983), .B2(new_n977), .ZN(G1352gat));
  OR3_X1    g783(.A1(new_n980), .A2(G204gat), .A3(new_n661), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n987), .B1(new_n976), .B2(new_n661), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n975), .A2(KEYINPUT126), .A3(new_n660), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n988), .A2(G204gat), .A3(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n985), .A2(KEYINPUT62), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n986), .A2(new_n990), .A3(new_n991), .ZN(G1353gat));
  NOR2_X1   g791(.A1(new_n581), .A2(G211gat), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n981), .A2(new_n982), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n975), .A2(new_n689), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n995), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n996));
  INV_X1    g795(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g796(.A(KEYINPUT63), .B1(new_n995), .B2(G211gat), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n994), .B1(new_n997), .B2(new_n998), .ZN(G1354gat));
  NAND3_X1  g798(.A1(new_n981), .A2(new_n624), .A3(new_n982), .ZN(new_n1000));
  INV_X1    g799(.A(G218gat), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n624), .A2(G218gat), .ZN(new_n1002));
  XNOR2_X1  g801(.A(new_n1002), .B(KEYINPUT127), .ZN(new_n1003));
  AOI22_X1  g802(.A1(new_n1000), .A2(new_n1001), .B1(new_n975), .B2(new_n1003), .ZN(G1355gat));
endmodule


