//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n733, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n811, new_n812, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n898,
    new_n899, new_n901, new_n902, new_n903, new_n904, new_n905, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935;
  INV_X1    g000(.A(KEYINPUT1), .ZN(new_n202));
  OAI21_X1  g001(.A(new_n202), .B1(G113gat), .B2(G120gat), .ZN(new_n203));
  AOI21_X1  g002(.A(new_n203), .B1(G113gat), .B2(G120gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(KEYINPUT74), .ZN(new_n205));
  INV_X1    g004(.A(G127gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(G134gat), .ZN(new_n207));
  INV_X1    g006(.A(G134gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G127gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n205), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n204), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(G127gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n206), .A2(G134gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G113gat), .ZN(new_n215));
  INV_X1    g014(.A(G120gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n214), .B(new_n205), .C1(new_n217), .C2(new_n203), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(G169gat), .ZN(new_n220));
  INV_X1    g019(.A(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(KEYINPUT26), .ZN(new_n223));
  AND2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n222), .A2(KEYINPUT26), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n225), .A2(new_n226), .B1(G183gat), .B2(G190gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT28), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT27), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT71), .B1(new_n229), .B2(G183gat), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT71), .ZN(new_n231));
  INV_X1    g030(.A(G183gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n232), .A3(KEYINPUT27), .ZN(new_n233));
  INV_X1    g032(.A(G190gat), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  OR2_X1    g034(.A1(KEYINPUT72), .A2(KEYINPUT27), .ZN(new_n236));
  NAND2_X1  g035(.A1(KEYINPUT72), .A2(KEYINPUT27), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n232), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n228), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT73), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT27), .B(G183gat), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n241), .A2(KEYINPUT28), .A3(new_n234), .ZN(new_n242));
  AND3_X1   g041(.A1(new_n239), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n240), .B1(new_n239), .B2(new_n242), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n227), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT23), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n224), .B1(new_n222), .B2(new_n246), .ZN(new_n247));
  OAI211_X1 g046(.A(new_n247), .B(KEYINPUT25), .C1(new_n246), .C2(new_n222), .ZN(new_n248));
  NAND3_X1  g047(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252));
  NOR3_X1   g051(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n248), .A2(new_n253), .ZN(new_n254));
  OR2_X1    g053(.A1(KEYINPUT68), .A2(G176gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(KEYINPUT68), .A2(G176gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(KEYINPUT23), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n220), .A2(KEYINPUT67), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT67), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G169gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n247), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n247), .B(KEYINPUT69), .C1(new_n257), .C2(new_n261), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n252), .A2(KEYINPUT66), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT66), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n267), .B1(G183gat), .B2(G190gat), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n251), .A2(KEYINPUT65), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n249), .A2(KEYINPUT64), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n273), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G183gat), .A2(G190gat), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT24), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n276), .A2(KEYINPUT65), .A3(new_n277), .ZN(new_n278));
  NAND4_X1  g077(.A1(new_n269), .A2(new_n271), .A3(new_n275), .A4(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n265), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT25), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n254), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n245), .B1(new_n282), .B2(KEYINPUT70), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT70), .ZN(new_n284));
  AOI211_X1 g083(.A(new_n284), .B(new_n254), .C1(new_n280), .C2(new_n281), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n219), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n266), .A2(new_n278), .A3(new_n268), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n287), .A2(new_n270), .ZN(new_n288));
  AOI22_X1  g087(.A1(new_n288), .A2(new_n275), .B1(new_n262), .B2(new_n263), .ZN(new_n289));
  AOI21_X1  g088(.A(KEYINPUT25), .B1(new_n289), .B2(new_n265), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n284), .B1(new_n290), .B2(new_n254), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n282), .A2(KEYINPUT70), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n211), .A2(new_n218), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .A4(new_n245), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n286), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G227gat), .A2(G233gat), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(KEYINPUT32), .ZN(new_n299));
  XOR2_X1   g098(.A(KEYINPUT75), .B(KEYINPUT33), .Z(new_n300));
  NAND2_X1  g099(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G15gat), .B(G43gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(G71gat), .B(G99gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n302), .B(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n299), .A2(new_n301), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n286), .A2(new_n296), .A3(new_n294), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT76), .B1(new_n307), .B2(KEYINPUT34), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(KEYINPUT34), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n298), .B(KEYINPUT32), .C1(new_n304), .C2(new_n300), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n307), .A2(KEYINPUT76), .A3(KEYINPUT34), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n306), .A2(new_n310), .A3(new_n311), .A4(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT77), .ZN(new_n314));
  INV_X1    g113(.A(new_n312), .ZN(new_n315));
  NOR3_X1   g114(.A1(new_n315), .A2(new_n309), .A3(new_n308), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT77), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n316), .A2(new_n317), .A3(new_n311), .A4(new_n306), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n306), .A2(new_n311), .ZN(new_n320));
  OR2_X1    g119(.A1(new_n320), .A2(new_n316), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT80), .ZN(new_n322));
  INV_X1    g121(.A(G141gat), .ZN(new_n323));
  INV_X1    g122(.A(G148gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(G141gat), .A2(G148gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n328), .B1(G155gat), .B2(G162gat), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n322), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G155gat), .B(G162gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n322), .B(new_n331), .C1(new_n327), .C2(new_n329), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  XNOR2_X1  g134(.A(G197gat), .B(G204gat), .ZN(new_n336));
  INV_X1    g135(.A(G211gat), .ZN(new_n337));
  INV_X1    g136(.A(G218gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n336), .B1(KEYINPUT22), .B2(new_n339), .ZN(new_n340));
  XOR2_X1   g139(.A(G211gat), .B(G218gat), .Z(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT29), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT3), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n335), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n335), .A2(new_n345), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n342), .B1(new_n347), .B2(new_n343), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(G50gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(G78gat), .B(G106gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT31), .ZN(new_n352));
  NAND2_X1  g151(.A1(G228gat), .A2(G233gat), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n353), .B(G22gat), .Z(new_n354));
  XNOR2_X1  g153(.A(new_n352), .B(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n350), .A2(new_n355), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n319), .A2(new_n321), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n293), .A2(new_n335), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT4), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT4), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n293), .A2(new_n335), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT5), .ZN(new_n365));
  NAND2_X1  g164(.A1(G225gat), .A2(G233gat), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT81), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n219), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n333), .A2(KEYINPUT3), .A3(new_n334), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n211), .A2(new_n218), .A3(KEYINPUT81), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n347), .A2(new_n368), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n364), .A2(new_n365), .A3(new_n366), .A4(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n361), .A2(new_n363), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n360), .A2(KEYINPUT82), .A3(KEYINPUT4), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n366), .A4(new_n371), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n368), .A2(new_n370), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n360), .B1(new_n378), .B2(new_n335), .ZN(new_n379));
  INV_X1    g178(.A(new_n366), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n365), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT83), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n377), .A2(KEYINPUT83), .A3(new_n381), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n373), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT0), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n388), .B(G57gat), .ZN(new_n389));
  INV_X1    g188(.A(G85gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(KEYINPUT6), .B1(new_n386), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n392), .B1(new_n391), .B2(new_n386), .ZN(new_n393));
  INV_X1    g192(.A(new_n385), .ZN(new_n394));
  AOI21_X1  g193(.A(KEYINPUT83), .B1(new_n377), .B2(new_n381), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n372), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n391), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(KEYINPUT6), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(G8gat), .B(G36gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n400), .B(G64gat), .ZN(new_n401));
  INV_X1    g200(.A(G92gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(new_n401), .B(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n282), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n245), .ZN(new_n405));
  NAND2_X1  g204(.A1(G226gat), .A2(G233gat), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n343), .B1(new_n283), .B2(new_n285), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(new_n406), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n409), .B1(new_n411), .B2(KEYINPUT79), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n291), .A2(new_n292), .A3(new_n245), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n407), .B1(new_n413), .B2(new_n343), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n342), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n342), .ZN(new_n418));
  OR2_X1    g217(.A1(new_n413), .A2(new_n406), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n405), .A2(new_n343), .A3(new_n406), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(KEYINPUT30), .B(new_n403), .C1(new_n417), .C2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n408), .B1(new_n414), .B2(new_n415), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n411), .A2(KEYINPUT79), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n418), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n403), .A2(KEYINPUT30), .ZN(new_n426));
  OR2_X1    g225(.A1(new_n403), .A2(KEYINPUT30), .ZN(new_n427));
  INV_X1    g226(.A(new_n421), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n422), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n399), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT35), .B1(new_n359), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n396), .A2(KEYINPUT86), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT86), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n386), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n391), .B1(new_n433), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n392), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT88), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n384), .A2(new_n385), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n434), .B1(new_n439), .B2(new_n372), .ZN(new_n440));
  AOI211_X1 g239(.A(KEYINPUT86), .B(new_n373), .C1(new_n384), .C2(new_n385), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n397), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT88), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(new_n443), .A3(new_n392), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n438), .A2(new_n444), .A3(new_n398), .ZN(new_n445));
  INV_X1    g244(.A(new_n358), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT90), .B(KEYINPUT35), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT84), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n422), .A2(new_n429), .A3(KEYINPUT84), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  OAI211_X1 g252(.A(new_n445), .B(new_n448), .C1(new_n451), .C2(new_n453), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n314), .A2(KEYINPUT78), .A3(new_n318), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT78), .B1(new_n314), .B2(new_n318), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n321), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n432), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT87), .ZN(new_n459));
  OR2_X1    g258(.A1(new_n379), .A2(new_n380), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT85), .B1(new_n460), .B2(KEYINPUT39), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n366), .B1(new_n364), .B2(new_n371), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(KEYINPUT85), .A3(KEYINPUT39), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT39), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g266(.A1(new_n465), .A2(KEYINPUT40), .A3(new_n391), .A4(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  INV_X1    g268(.A(new_n464), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n470), .A2(new_n461), .A3(new_n462), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n467), .A2(new_n391), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n468), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n474), .A2(new_n436), .ZN(new_n475));
  NAND4_X1  g274(.A1(new_n450), .A2(new_n459), .A3(new_n452), .A4(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n450), .A2(new_n452), .A3(new_n475), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT87), .ZN(new_n478));
  INV_X1    g277(.A(new_n398), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n442), .A2(new_n392), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n480), .B2(KEYINPUT88), .ZN(new_n481));
  XOR2_X1   g280(.A(KEYINPUT89), .B(KEYINPUT37), .Z(new_n482));
  NOR3_X1   g281(.A1(new_n417), .A2(new_n421), .A3(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT37), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n425), .B2(new_n428), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT38), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  OR3_X1    g285(.A1(new_n417), .A2(new_n421), .A3(new_n482), .ZN(new_n487));
  OR2_X1    g286(.A1(new_n403), .A2(KEYINPUT38), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n342), .B1(new_n423), .B2(new_n424), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n419), .A2(new_n420), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n484), .B1(new_n490), .B2(new_n418), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n488), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT38), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(new_n417), .B2(new_n421), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n487), .A2(new_n492), .B1(new_n494), .B2(new_n403), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n481), .A2(new_n486), .A3(new_n444), .A4(new_n495), .ZN(new_n496));
  AND4_X1   g295(.A1(new_n476), .A2(new_n478), .A3(new_n358), .A4(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n498), .B(new_n321), .C1(new_n455), .C2(new_n456), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n319), .A2(new_n321), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT36), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n431), .A2(new_n446), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n499), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n458), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT91), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n458), .B(KEYINPUT91), .C1(new_n497), .C2(new_n503), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G15gat), .B(G22gat), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT96), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT16), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(G1gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  NOR3_X1   g312(.A1(new_n510), .A2(new_n511), .A3(G1gat), .ZN(new_n514));
  OAI22_X1  g313(.A1(new_n513), .A2(new_n514), .B1(G1gat), .B2(new_n509), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT97), .B1(new_n509), .B2(G1gat), .ZN(new_n516));
  INV_X1    g315(.A(G8gat), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n515), .B(new_n518), .ZN(new_n519));
  XOR2_X1   g318(.A(G43gat), .B(G50gat), .Z(new_n520));
  INV_X1    g319(.A(KEYINPUT15), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT94), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n520), .A2(new_n521), .ZN(new_n524));
  INV_X1    g323(.A(G29gat), .ZN(new_n525));
  INV_X1    g324(.A(G36gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT14), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT14), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n527), .B(new_n529), .C1(new_n525), .C2(new_n526), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n523), .A2(new_n524), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n530), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT93), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT95), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(KEYINPUT17), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n538), .B1(new_n534), .B2(new_n535), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n519), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT98), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT98), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G229gat), .A2(G233gat), .ZN(new_n545));
  XOR2_X1   g344(.A(new_n545), .B(KEYINPUT99), .Z(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n519), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n534), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n542), .A2(new_n544), .A3(new_n547), .A4(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT18), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n550), .B1(new_n540), .B2(new_n543), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n555), .A2(KEYINPUT18), .A3(new_n547), .A4(new_n544), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n534), .B(new_n519), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n546), .B(KEYINPUT13), .Z(new_n558));
  OR2_X1    g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n553), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n561));
  XNOR2_X1  g360(.A(G113gat), .B(G141gat), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(KEYINPUT11), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(new_n220), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(G197gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT12), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n560), .A2(new_n561), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n567), .B1(new_n560), .B2(new_n561), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G190gat), .B(G218gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n537), .A2(new_n539), .ZN(new_n572));
  NAND2_X1  g371(.A1(G99gat), .A2(G106gat), .ZN(new_n573));
  AOI22_X1  g372(.A1(KEYINPUT8), .A2(new_n573), .B1(new_n390), .B2(new_n402), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT104), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G85gat), .A2(G92gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(KEYINPUT7), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G99gat), .B(G106gat), .Z(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT105), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n579), .A2(new_n580), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n572), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n571), .A2(KEYINPUT106), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT41), .ZN(new_n587));
  NAND2_X1  g386(.A1(G232gat), .A2(G233gat), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n584), .ZN(new_n590));
  INV_X1    g389(.A(new_n534), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI211_X1 g391(.A(KEYINPUT106), .B(new_n571), .C1(new_n585), .C2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n585), .A2(new_n592), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n571), .A2(KEYINPUT106), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n588), .A2(new_n587), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT103), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(new_n208), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(G162gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n601), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n603), .B1(new_n593), .B2(new_n596), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(KEYINPUT100), .B(G57gat), .Z(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(G64gat), .ZN(new_n608));
  INV_X1    g407(.A(G57gat), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n608), .B1(new_n609), .B2(G64gat), .ZN(new_n610));
  AND2_X1   g409(.A1(G71gat), .A2(G78gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n611), .A2(KEYINPUT9), .ZN(new_n612));
  NOR2_X1   g411(.A1(G71gat), .A2(G78gat), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n612), .B1(new_n615), .B2(KEYINPUT101), .ZN(new_n616));
  OAI211_X1 g415(.A(new_n610), .B(new_n616), .C1(KEYINPUT101), .C2(new_n615), .ZN(new_n617));
  XNOR2_X1  g416(.A(G57gat), .B(G64gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT9), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n614), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT21), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g424(.A(G127gat), .B(G155gat), .Z(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT20), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n625), .B(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n548), .B1(new_n621), .B2(new_n622), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G183gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n628), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT102), .B(KEYINPUT19), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(G211gat), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n631), .A2(new_n633), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n584), .A2(new_n621), .ZN(new_n637));
  INV_X1    g436(.A(new_n621), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(new_n583), .A3(new_n581), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT107), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT10), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n637), .A2(new_n645), .A3(new_n639), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n590), .A2(KEYINPUT10), .A3(new_n638), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n641), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(G148gat), .ZN(new_n651));
  XOR2_X1   g450(.A(KEYINPUT108), .B(G120gat), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n644), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n649), .A2(new_n643), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n653), .B(KEYINPUT109), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n606), .A2(new_n636), .A3(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n570), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n508), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n399), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g464(.A1(new_n451), .A2(new_n453), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT16), .B(G8gat), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT42), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n667), .A2(G8gat), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n669), .A2(new_n670), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(G1325gat));
  INV_X1    g473(.A(new_n457), .ZN(new_n675));
  AOI21_X1  g474(.A(G15gat), .B1(new_n662), .B2(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(KEYINPUT110), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n499), .A2(new_n501), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n679), .A2(G15gat), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n677), .B1(new_n662), .B2(new_n680), .ZN(G1326gat));
  NAND2_X1  g480(.A1(new_n662), .A2(new_n446), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT43), .B(G22gat), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(G1327gat));
  NOR3_X1   g483(.A1(new_n570), .A2(new_n636), .A3(new_n658), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n508), .A2(new_n605), .A3(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n686), .A2(G29gat), .A3(new_n399), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n504), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT113), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n605), .B(new_n691), .ZN(new_n692));
  OR3_X1    g491(.A1(new_n690), .A2(KEYINPUT44), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n506), .A2(new_n507), .A3(new_n605), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n694), .A2(KEYINPUT112), .A3(KEYINPUT44), .ZN(new_n695));
  AOI21_X1  g494(.A(KEYINPUT112), .B1(new_n694), .B2(KEYINPUT44), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n697), .A2(new_n685), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n698), .A2(new_n663), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n689), .B1(new_n699), .B2(new_n525), .ZN(G1328gat));
  INV_X1    g499(.A(new_n666), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n686), .A2(G36gat), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT46), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n698), .A2(new_n666), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(new_n526), .ZN(G1329gat));
  OR2_X1    g504(.A1(new_n457), .A2(G43gat), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n686), .A2(new_n706), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n697), .A2(new_n679), .A3(new_n685), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(new_n708), .B2(G43gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g509(.A1(new_n358), .A2(G50gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(KEYINPUT114), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n686), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n697), .A2(new_n446), .A3(new_n685), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n714), .B2(G50gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT48), .ZN(G1331gat));
  AND3_X1   g515(.A1(new_n553), .A2(new_n556), .A3(new_n559), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n566), .B1(new_n717), .B2(KEYINPUT92), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n560), .A2(new_n561), .A3(new_n567), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n606), .A2(new_n636), .A3(new_n658), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n690), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n663), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(new_n607), .Z(G1332gat));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n666), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n725), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n726));
  XOR2_X1   g525(.A(KEYINPUT49), .B(G64gat), .Z(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n725), .B2(new_n727), .ZN(G1333gat));
  NAND2_X1  g527(.A1(new_n722), .A2(new_n679), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n457), .A2(G71gat), .ZN(new_n730));
  AOI22_X1  g529(.A1(new_n729), .A2(G71gat), .B1(new_n722), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g531(.A1(new_n722), .A2(new_n446), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(G78gat), .ZN(G1335gat));
  INV_X1    g533(.A(new_n636), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n570), .A2(new_n735), .A3(new_n605), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n690), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g536(.A1(new_n737), .A2(KEYINPUT51), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(KEYINPUT51), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n659), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n740), .A2(new_n390), .A3(new_n663), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n720), .A2(new_n636), .A3(new_n659), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n697), .A2(new_n742), .ZN(new_n743));
  AND2_X1   g542(.A1(new_n743), .A2(new_n663), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n741), .B1(new_n744), .B2(new_n390), .ZN(G1336gat));
  NOR2_X1   g544(.A1(new_n701), .A2(G92gat), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  AOI211_X1 g546(.A(new_n659), .B(new_n747), .C1(new_n738), .C2(new_n739), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n697), .A2(new_n666), .A3(new_n742), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n748), .B1(new_n749), .B2(G92gat), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT115), .ZN(new_n751));
  AND3_X1   g550(.A1(new_n750), .A2(new_n751), .A3(KEYINPUT52), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(KEYINPUT52), .ZN(new_n753));
  AND2_X1   g552(.A1(new_n751), .A2(KEYINPUT52), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n750), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n752), .A2(new_n755), .ZN(G1337gat));
  AOI21_X1  g555(.A(G99gat), .B1(new_n740), .B2(new_n675), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n679), .A2(G99gat), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n757), .B1(new_n743), .B2(new_n758), .ZN(G1338gat));
  NAND3_X1  g558(.A1(new_n697), .A2(new_n446), .A3(new_n742), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G106gat), .ZN(new_n761));
  INV_X1    g560(.A(G106gat), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n740), .A2(new_n762), .A3(new_n446), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT116), .B(KEYINPUT53), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1339gat));
  NOR2_X1   g565(.A1(new_n720), .A2(new_n660), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n544), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n546), .B1(new_n769), .B2(new_n554), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT117), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT117), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n772), .B(new_n546), .C1(new_n769), .C2(new_n554), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n557), .A2(new_n558), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  AOI22_X1  g574(.A1(new_n717), .A2(new_n566), .B1(new_n775), .B2(new_n565), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n658), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n646), .A2(new_n642), .A3(new_n647), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n649), .A2(KEYINPUT54), .A3(new_n778), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n642), .B1(new_n646), .B2(new_n647), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT54), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n653), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n779), .A2(KEYINPUT55), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n654), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n779), .A2(new_n782), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n784), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n777), .B1(new_n570), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n692), .ZN(new_n790));
  INV_X1    g589(.A(new_n692), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(new_n776), .A3(new_n787), .ZN(new_n792));
  AND2_X1   g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n768), .B1(new_n793), .B2(new_n636), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n358), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n795), .A2(KEYINPUT118), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(KEYINPUT118), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n798), .A2(new_n663), .A3(new_n701), .A4(new_n675), .ZN(new_n799));
  OAI21_X1  g598(.A(G113gat), .B1(new_n799), .B2(new_n570), .ZN(new_n800));
  AND2_X1   g599(.A1(new_n794), .A2(new_n663), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n666), .A2(new_n359), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n570), .A2(G113gat), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n804), .B(KEYINPUT119), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n800), .B1(new_n803), .B2(new_n805), .ZN(G1340gat));
  NOR3_X1   g605(.A1(new_n799), .A2(new_n216), .A3(new_n659), .ZN(new_n807));
  INV_X1    g606(.A(new_n803), .ZN(new_n808));
  AOI21_X1  g607(.A(G120gat), .B1(new_n808), .B2(new_n658), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n807), .A2(new_n809), .ZN(G1341gat));
  OAI21_X1  g609(.A(G127gat), .B1(new_n799), .B2(new_n735), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n808), .A2(new_n206), .A3(new_n636), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1342gat));
  NOR3_X1   g612(.A1(new_n803), .A2(G134gat), .A3(new_n606), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT56), .ZN(new_n815));
  OAI21_X1  g614(.A(G134gat), .B1(new_n799), .B2(new_n606), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(G1343gat));
  NOR2_X1   g616(.A1(new_n666), .A2(new_n358), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n801), .A2(new_n678), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n820), .A2(new_n323), .A3(new_n720), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n794), .A2(new_n822), .A3(new_n446), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n679), .A2(new_n399), .A3(new_n666), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n786), .A2(new_n785), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT120), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n654), .A2(new_n783), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n786), .A2(new_n829), .A3(new_n785), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n831), .B1(new_n568), .B2(new_n569), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n605), .B1(new_n832), .B2(new_n777), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n834), .A2(new_n792), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n768), .B1(new_n835), .B2(new_n636), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n822), .B1(new_n836), .B2(new_n446), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n825), .A2(new_n837), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n838), .A2(new_n570), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n821), .B1(new_n839), .B2(new_n323), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(KEYINPUT58), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n842), .B(new_n821), .C1(new_n839), .C2(new_n323), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(G1344gat));
  NOR3_X1   g643(.A1(new_n819), .A2(G148gat), .A3(new_n659), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT121), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT59), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n794), .A2(new_n446), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT57), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT124), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT123), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n787), .A2(new_n851), .A3(new_n605), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n605), .A2(new_n828), .A3(new_n826), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT123), .ZN(new_n854));
  AND3_X1   g653(.A1(new_n852), .A2(new_n854), .A3(new_n776), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n850), .B1(new_n833), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(new_n854), .A3(new_n776), .ZN(new_n857));
  AOI22_X1  g656(.A1(new_n720), .A2(new_n831), .B1(new_n776), .B2(new_n658), .ZN(new_n858));
  OAI211_X1 g657(.A(KEYINPUT124), .B(new_n857), .C1(new_n858), .C2(new_n605), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n856), .A2(new_n735), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(new_n768), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n446), .ZN(new_n862));
  AOI21_X1  g661(.A(KEYINPUT125), .B1(new_n862), .B2(new_n822), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n358), .B1(new_n860), .B2(new_n768), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT125), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT57), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n849), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n658), .A3(new_n824), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n847), .B1(new_n868), .B2(G148gat), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n324), .A2(KEYINPUT59), .ZN(new_n870));
  OAI211_X1 g669(.A(KEYINPUT122), .B(new_n870), .C1(new_n838), .C2(new_n659), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n825), .A2(new_n837), .A3(new_n659), .ZN(new_n873));
  INV_X1    g672(.A(new_n870), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n846), .B1(new_n869), .B2(new_n876), .ZN(G1345gat));
  OAI21_X1  g676(.A(G155gat), .B1(new_n838), .B2(new_n735), .ZN(new_n878));
  OR3_X1    g677(.A1(new_n819), .A2(G155gat), .A3(new_n735), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1346gat));
  OAI21_X1  g679(.A(G162gat), .B1(new_n838), .B2(new_n692), .ZN(new_n881));
  OR3_X1    g680(.A1(new_n819), .A2(G162gat), .A3(new_n606), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(G1347gat));
  NOR2_X1   g682(.A1(new_n701), .A2(new_n663), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n359), .ZN(new_n886));
  AND2_X1   g685(.A1(new_n794), .A2(new_n886), .ZN(new_n887));
  XOR2_X1   g686(.A(new_n887), .B(KEYINPUT126), .Z(new_n888));
  NAND4_X1  g687(.A1(new_n888), .A2(new_n258), .A3(new_n260), .A4(new_n720), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT127), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n885), .A2(new_n457), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n892), .B1(new_n796), .B2(new_n797), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n720), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n890), .B1(new_n894), .B2(G169gat), .ZN(new_n895));
  AOI211_X1 g694(.A(KEYINPUT127), .B(new_n220), .C1(new_n893), .C2(new_n720), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n889), .B1(new_n895), .B2(new_n896), .ZN(G1348gat));
  AOI21_X1  g696(.A(G176gat), .B1(new_n888), .B2(new_n658), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n659), .B1(new_n255), .B2(new_n256), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n898), .B1(new_n893), .B2(new_n899), .ZN(G1349gat));
  AOI21_X1  g699(.A(new_n232), .B1(new_n893), .B2(new_n636), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n887), .A2(new_n241), .A3(new_n636), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  OR3_X1    g702(.A1(new_n901), .A2(KEYINPUT60), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT60), .B1(new_n901), .B2(new_n903), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(G1350gat));
  NAND3_X1  g705(.A1(new_n888), .A2(new_n234), .A3(new_n791), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n605), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(G190gat), .ZN(new_n910));
  AOI211_X1 g709(.A(KEYINPUT61), .B(new_n234), .C1(new_n893), .C2(new_n605), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(G1351gat));
  NOR2_X1   g711(.A1(new_n679), .A2(new_n885), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n848), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(G197gat), .B1(new_n914), .B2(new_n720), .ZN(new_n915));
  INV_X1    g714(.A(new_n913), .ZN(new_n916));
  INV_X1    g715(.A(new_n866), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n865), .B1(new_n864), .B2(KEYINPUT57), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n916), .B1(new_n919), .B2(new_n849), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n720), .A2(G197gat), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n915), .B1(new_n920), .B2(new_n921), .ZN(G1352gat));
  INV_X1    g721(.A(G204gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n914), .A2(new_n923), .A3(new_n658), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT62), .ZN(new_n925));
  OR2_X1    g724(.A1(new_n924), .A2(KEYINPUT62), .ZN(new_n926));
  AND3_X1   g725(.A1(new_n867), .A2(new_n658), .A3(new_n913), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n925), .B(new_n926), .C1(new_n927), .C2(new_n923), .ZN(G1353gat));
  NAND3_X1  g727(.A1(new_n914), .A2(new_n337), .A3(new_n636), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n867), .A2(new_n636), .A3(new_n913), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT63), .B1(new_n930), .B2(G211gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1354gat));
  AOI21_X1  g732(.A(G218gat), .B1(new_n914), .B2(new_n791), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n606), .A2(new_n338), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n934), .B1(new_n920), .B2(new_n935), .ZN(G1355gat));
endmodule


