

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U555 ( .A(n982), .ZN(n764) );
  NAND2_X1 U556 ( .A1(n523), .A2(n767), .ZN(n773) );
  INV_X1 U557 ( .A(n995), .ZN(n771) );
  NOR2_X1 U558 ( .A1(G651), .A2(G543), .ZN(n659) );
  AND2_X1 U559 ( .A1(n772), .A2(n771), .ZN(n521) );
  XOR2_X1 U560 ( .A(KEYINPUT14), .B(n577), .Z(n522) );
  NAND2_X1 U561 ( .A1(n766), .A2(n765), .ZN(n523) );
  INV_X1 U562 ( .A(KEYINPUT29), .ZN(n727) );
  NAND2_X1 U563 ( .A1(n747), .A2(n746), .ZN(n757) );
  NOR2_X1 U564 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U565 ( .A1(G651), .A2(n638), .ZN(n656) );
  NOR2_X2 U566 ( .A1(G2105), .A2(n546), .ZN(n906) );
  XOR2_X1 U567 ( .A(KEYINPUT1), .B(n530), .Z(n662) );
  AND2_X1 U568 ( .A1(n550), .A2(n549), .ZN(G160) );
  XOR2_X1 U569 ( .A(G543), .B(KEYINPUT0), .Z(n638) );
  INV_X1 U570 ( .A(G651), .ZN(n529) );
  NOR2_X1 U571 ( .A1(n638), .A2(n529), .ZN(n658) );
  NAND2_X1 U572 ( .A1(n658), .A2(G76), .ZN(n524) );
  XNOR2_X1 U573 ( .A(KEYINPUT76), .B(n524), .ZN(n527) );
  NAND2_X1 U574 ( .A1(n659), .A2(G89), .ZN(n525) );
  XNOR2_X1 U575 ( .A(KEYINPUT4), .B(n525), .ZN(n526) );
  NAND2_X1 U576 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U577 ( .A(n528), .B(KEYINPUT5), .ZN(n535) );
  NAND2_X1 U578 ( .A1(G51), .A2(n656), .ZN(n532) );
  NOR2_X1 U579 ( .A1(G543), .A2(n529), .ZN(n530) );
  NAND2_X1 U580 ( .A1(G63), .A2(n662), .ZN(n531) );
  NAND2_X1 U581 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U582 ( .A(KEYINPUT6), .B(n533), .Z(n534) );
  NAND2_X1 U583 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U584 ( .A(n536), .B(KEYINPUT7), .ZN(G168) );
  XNOR2_X1 U585 ( .A(G168), .B(KEYINPUT8), .ZN(n537) );
  XNOR2_X1 U586 ( .A(n537), .B(KEYINPUT77), .ZN(G286) );
  INV_X1 U587 ( .A(G2104), .ZN(n546) );
  NAND2_X1 U588 ( .A1(G101), .A2(n906), .ZN(n538) );
  XOR2_X1 U589 ( .A(KEYINPUT23), .B(n538), .Z(n550) );
  NOR2_X1 U590 ( .A1(G2105), .A2(G2104), .ZN(n539) );
  XNOR2_X1 U591 ( .A(n539), .B(KEYINPUT66), .ZN(n541) );
  XNOR2_X1 U592 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n540) );
  XNOR2_X1 U593 ( .A(n541), .B(n540), .ZN(n567) );
  NAND2_X1 U594 ( .A1(G137), .A2(n567), .ZN(n543) );
  AND2_X1 U595 ( .A1(G2105), .A2(G2104), .ZN(n903) );
  NAND2_X1 U596 ( .A1(G113), .A2(n903), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(n545) );
  INV_X1 U598 ( .A(KEYINPUT68), .ZN(n544) );
  XNOR2_X1 U599 ( .A(n545), .B(n544), .ZN(n548) );
  AND2_X1 U600 ( .A1(n546), .A2(G2105), .ZN(n902) );
  NAND2_X1 U601 ( .A1(n902), .A2(G125), .ZN(n547) );
  AND2_X1 U602 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U603 ( .A(G2443), .B(G2446), .Z(n552) );
  XNOR2_X1 U604 ( .A(G2427), .B(G2451), .ZN(n551) );
  XNOR2_X1 U605 ( .A(n552), .B(n551), .ZN(n558) );
  XOR2_X1 U606 ( .A(G2430), .B(G2454), .Z(n554) );
  XNOR2_X1 U607 ( .A(G1348), .B(G1341), .ZN(n553) );
  XNOR2_X1 U608 ( .A(n554), .B(n553), .ZN(n556) );
  XOR2_X1 U609 ( .A(G2435), .B(G2438), .Z(n555) );
  XNOR2_X1 U610 ( .A(n556), .B(n555), .ZN(n557) );
  XOR2_X1 U611 ( .A(n558), .B(n557), .Z(n559) );
  AND2_X1 U612 ( .A1(G14), .A2(n559), .ZN(G401) );
  AND2_X1 U613 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U614 ( .A(G57), .ZN(G237) );
  NAND2_X1 U615 ( .A1(G52), .A2(n656), .ZN(n561) );
  NAND2_X1 U616 ( .A1(G64), .A2(n662), .ZN(n560) );
  NAND2_X1 U617 ( .A1(n561), .A2(n560), .ZN(n566) );
  NAND2_X1 U618 ( .A1(G77), .A2(n658), .ZN(n563) );
  NAND2_X1 U619 ( .A1(G90), .A2(n659), .ZN(n562) );
  NAND2_X1 U620 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U621 ( .A(KEYINPUT9), .B(n564), .Z(n565) );
  NOR2_X1 U622 ( .A1(n566), .A2(n565), .ZN(G171) );
  NAND2_X1 U623 ( .A1(n906), .A2(G102), .ZN(n569) );
  BUF_X1 U624 ( .A(n567), .Z(n613) );
  NAND2_X1 U625 ( .A1(G138), .A2(n613), .ZN(n568) );
  NAND2_X1 U626 ( .A1(n569), .A2(n568), .ZN(n573) );
  NAND2_X1 U627 ( .A1(G126), .A2(n902), .ZN(n571) );
  NAND2_X1 U628 ( .A1(G114), .A2(n903), .ZN(n570) );
  NAND2_X1 U629 ( .A1(n571), .A2(n570), .ZN(n572) );
  NOR2_X1 U630 ( .A1(n573), .A2(n572), .ZN(G164) );
  NAND2_X1 U631 ( .A1(G7), .A2(G661), .ZN(n574) );
  XNOR2_X1 U632 ( .A(n574), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U633 ( .A(G223), .ZN(n843) );
  NAND2_X1 U634 ( .A1(n843), .A2(G567), .ZN(n575) );
  XNOR2_X1 U635 ( .A(n575), .B(KEYINPUT71), .ZN(n576) );
  XNOR2_X1 U636 ( .A(KEYINPUT11), .B(n576), .ZN(G234) );
  NAND2_X1 U637 ( .A1(G56), .A2(n662), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n659), .A2(G81), .ZN(n578) );
  XNOR2_X1 U639 ( .A(n578), .B(KEYINPUT12), .ZN(n580) );
  NAND2_X1 U640 ( .A1(G68), .A2(n658), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U642 ( .A(KEYINPUT13), .B(n581), .Z(n582) );
  NOR2_X1 U643 ( .A1(n522), .A2(n582), .ZN(n584) );
  NAND2_X1 U644 ( .A1(n656), .A2(G43), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n584), .A2(n583), .ZN(n979) );
  INV_X1 U646 ( .A(G860), .ZN(n627) );
  NOR2_X1 U647 ( .A1(n979), .A2(n627), .ZN(n585) );
  XOR2_X1 U648 ( .A(KEYINPUT72), .B(n585), .Z(G153) );
  INV_X1 U649 ( .A(G868), .ZN(n604) );
  NOR2_X1 U650 ( .A1(n604), .A2(G171), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(KEYINPUT73), .ZN(n596) );
  NAND2_X1 U652 ( .A1(G92), .A2(n659), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G66), .A2(n662), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U655 ( .A1(G79), .A2(n658), .ZN(n590) );
  NAND2_X1 U656 ( .A1(G54), .A2(n656), .ZN(n589) );
  NAND2_X1 U657 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U658 ( .A1(n592), .A2(n591), .ZN(n594) );
  XNOR2_X1 U659 ( .A(KEYINPUT74), .B(KEYINPUT15), .ZN(n593) );
  XNOR2_X1 U660 ( .A(n594), .B(n593), .ZN(n849) );
  NAND2_X1 U661 ( .A1(n604), .A2(n849), .ZN(n595) );
  NAND2_X1 U662 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U663 ( .A(KEYINPUT75), .B(n597), .Z(G284) );
  NAND2_X1 U664 ( .A1(G53), .A2(n656), .ZN(n599) );
  NAND2_X1 U665 ( .A1(G65), .A2(n662), .ZN(n598) );
  NAND2_X1 U666 ( .A1(n599), .A2(n598), .ZN(n603) );
  NAND2_X1 U667 ( .A1(G78), .A2(n658), .ZN(n601) );
  NAND2_X1 U668 ( .A1(G91), .A2(n659), .ZN(n600) );
  NAND2_X1 U669 ( .A1(n601), .A2(n600), .ZN(n602) );
  NOR2_X1 U670 ( .A1(n603), .A2(n602), .ZN(n975) );
  INV_X1 U671 ( .A(n975), .ZN(G299) );
  NOR2_X1 U672 ( .A1(G286), .A2(n604), .ZN(n606) );
  NOR2_X1 U673 ( .A1(G868), .A2(G299), .ZN(n605) );
  NOR2_X1 U674 ( .A1(n606), .A2(n605), .ZN(G297) );
  NAND2_X1 U675 ( .A1(n627), .A2(G559), .ZN(n607) );
  INV_X1 U676 ( .A(n849), .ZN(n984) );
  NAND2_X1 U677 ( .A1(n607), .A2(n984), .ZN(n608) );
  XNOR2_X1 U678 ( .A(n608), .B(KEYINPUT16), .ZN(n609) );
  XNOR2_X1 U679 ( .A(KEYINPUT78), .B(n609), .ZN(G148) );
  NOR2_X1 U680 ( .A1(G868), .A2(n979), .ZN(n612) );
  NAND2_X1 U681 ( .A1(n984), .A2(G868), .ZN(n610) );
  NOR2_X1 U682 ( .A1(G559), .A2(n610), .ZN(n611) );
  NOR2_X1 U683 ( .A1(n612), .A2(n611), .ZN(G282) );
  NAND2_X1 U684 ( .A1(n613), .A2(G135), .ZN(n614) );
  XNOR2_X1 U685 ( .A(n614), .B(KEYINPUT80), .ZN(n618) );
  XOR2_X1 U686 ( .A(KEYINPUT79), .B(KEYINPUT18), .Z(n616) );
  NAND2_X1 U687 ( .A1(G123), .A2(n902), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n616), .B(n615), .ZN(n617) );
  NAND2_X1 U689 ( .A1(n618), .A2(n617), .ZN(n623) );
  NAND2_X1 U690 ( .A1(G111), .A2(n903), .ZN(n620) );
  NAND2_X1 U691 ( .A1(G99), .A2(n906), .ZN(n619) );
  NAND2_X1 U692 ( .A1(n620), .A2(n619), .ZN(n621) );
  XOR2_X1 U693 ( .A(KEYINPUT81), .B(n621), .Z(n622) );
  NOR2_X1 U694 ( .A1(n623), .A2(n622), .ZN(n933) );
  XOR2_X1 U695 ( .A(G2096), .B(n933), .Z(n624) );
  NOR2_X1 U696 ( .A1(G2100), .A2(n624), .ZN(n625) );
  XOR2_X1 U697 ( .A(KEYINPUT82), .B(n625), .Z(G156) );
  NAND2_X1 U698 ( .A1(n984), .A2(G559), .ZN(n626) );
  XOR2_X1 U699 ( .A(n979), .B(n626), .Z(n673) );
  NAND2_X1 U700 ( .A1(n627), .A2(n673), .ZN(n634) );
  NAND2_X1 U701 ( .A1(G55), .A2(n656), .ZN(n629) );
  NAND2_X1 U702 ( .A1(G67), .A2(n662), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n629), .A2(n628), .ZN(n633) );
  NAND2_X1 U704 ( .A1(G80), .A2(n658), .ZN(n631) );
  NAND2_X1 U705 ( .A1(G93), .A2(n659), .ZN(n630) );
  NAND2_X1 U706 ( .A1(n631), .A2(n630), .ZN(n632) );
  NOR2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n676) );
  XOR2_X1 U708 ( .A(n634), .B(n676), .Z(G145) );
  NAND2_X1 U709 ( .A1(G49), .A2(n656), .ZN(n636) );
  NAND2_X1 U710 ( .A1(G74), .A2(G651), .ZN(n635) );
  NAND2_X1 U711 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U712 ( .A1(n662), .A2(n637), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n638), .A2(G87), .ZN(n639) );
  NAND2_X1 U714 ( .A1(n640), .A2(n639), .ZN(G288) );
  NAND2_X1 U715 ( .A1(n658), .A2(G73), .ZN(n641) );
  XNOR2_X1 U716 ( .A(n641), .B(KEYINPUT2), .ZN(n648) );
  NAND2_X1 U717 ( .A1(G86), .A2(n659), .ZN(n643) );
  NAND2_X1 U718 ( .A1(G48), .A2(n656), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n646) );
  NAND2_X1 U720 ( .A1(G61), .A2(n662), .ZN(n644) );
  XNOR2_X1 U721 ( .A(KEYINPUT83), .B(n644), .ZN(n645) );
  NOR2_X1 U722 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(G305) );
  NAND2_X1 U724 ( .A1(G75), .A2(n658), .ZN(n650) );
  NAND2_X1 U725 ( .A1(G88), .A2(n659), .ZN(n649) );
  NAND2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n655) );
  NAND2_X1 U727 ( .A1(G62), .A2(n662), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n651), .B(KEYINPUT84), .ZN(n653) );
  NAND2_X1 U729 ( .A1(n656), .A2(G50), .ZN(n652) );
  NAND2_X1 U730 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U731 ( .A1(n655), .A2(n654), .ZN(G166) );
  INV_X1 U732 ( .A(G166), .ZN(G303) );
  NAND2_X1 U733 ( .A1(G47), .A2(n656), .ZN(n657) );
  XNOR2_X1 U734 ( .A(n657), .B(KEYINPUT70), .ZN(n667) );
  NAND2_X1 U735 ( .A1(G72), .A2(n658), .ZN(n661) );
  NAND2_X1 U736 ( .A1(G85), .A2(n659), .ZN(n660) );
  NAND2_X1 U737 ( .A1(n661), .A2(n660), .ZN(n665) );
  NAND2_X1 U738 ( .A1(G60), .A2(n662), .ZN(n663) );
  XNOR2_X1 U739 ( .A(KEYINPUT69), .B(n663), .ZN(n664) );
  NOR2_X1 U740 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U741 ( .A1(n667), .A2(n666), .ZN(G290) );
  XNOR2_X1 U742 ( .A(KEYINPUT19), .B(G288), .ZN(n672) );
  XNOR2_X1 U743 ( .A(n975), .B(n676), .ZN(n670) );
  XNOR2_X1 U744 ( .A(G305), .B(G303), .ZN(n668) );
  XNOR2_X1 U745 ( .A(n668), .B(G290), .ZN(n669) );
  XNOR2_X1 U746 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U747 ( .A(n672), .B(n671), .ZN(n852) );
  XNOR2_X1 U748 ( .A(n852), .B(n673), .ZN(n674) );
  NAND2_X1 U749 ( .A1(n674), .A2(G868), .ZN(n675) );
  XOR2_X1 U750 ( .A(KEYINPUT85), .B(n675), .Z(n678) );
  OR2_X1 U751 ( .A1(n676), .A2(G868), .ZN(n677) );
  NAND2_X1 U752 ( .A1(n678), .A2(n677), .ZN(G295) );
  NAND2_X1 U753 ( .A1(G2078), .A2(G2084), .ZN(n679) );
  XOR2_X1 U754 ( .A(KEYINPUT20), .B(n679), .Z(n680) );
  NAND2_X1 U755 ( .A1(G2090), .A2(n680), .ZN(n681) );
  XNOR2_X1 U756 ( .A(KEYINPUT21), .B(n681), .ZN(n682) );
  NAND2_X1 U757 ( .A1(n682), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U758 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U759 ( .A1(G132), .A2(G82), .ZN(n683) );
  XNOR2_X1 U760 ( .A(n683), .B(KEYINPUT22), .ZN(n684) );
  XNOR2_X1 U761 ( .A(n684), .B(KEYINPUT86), .ZN(n685) );
  NOR2_X1 U762 ( .A1(G218), .A2(n685), .ZN(n686) );
  NAND2_X1 U763 ( .A1(G96), .A2(n686), .ZN(n847) );
  NAND2_X1 U764 ( .A1(n847), .A2(G2106), .ZN(n690) );
  NAND2_X1 U765 ( .A1(G69), .A2(G120), .ZN(n687) );
  NOR2_X1 U766 ( .A1(G237), .A2(n687), .ZN(n688) );
  NAND2_X1 U767 ( .A1(G108), .A2(n688), .ZN(n848) );
  NAND2_X1 U768 ( .A1(n848), .A2(G567), .ZN(n689) );
  NAND2_X1 U769 ( .A1(n690), .A2(n689), .ZN(n925) );
  NAND2_X1 U770 ( .A1(G661), .A2(G483), .ZN(n691) );
  NOR2_X1 U771 ( .A1(n925), .A2(n691), .ZN(n846) );
  NAND2_X1 U772 ( .A1(n846), .A2(G36), .ZN(G176) );
  INV_X1 U773 ( .A(G171), .ZN(G301) );
  NOR2_X1 U774 ( .A1(G164), .A2(G1384), .ZN(n695) );
  NAND2_X1 U775 ( .A1(G160), .A2(G40), .ZN(n694) );
  NOR2_X1 U776 ( .A1(n695), .A2(n694), .ZN(n834) );
  XNOR2_X1 U777 ( .A(G1986), .B(G290), .ZN(n988) );
  NAND2_X1 U778 ( .A1(n834), .A2(n988), .ZN(n692) );
  XNOR2_X1 U779 ( .A(KEYINPUT87), .B(n692), .ZN(n788) );
  NOR2_X1 U780 ( .A1(G1976), .A2(G288), .ZN(n768) );
  NOR2_X1 U781 ( .A1(G1971), .A2(G303), .ZN(n693) );
  OR2_X1 U782 ( .A1(n768), .A2(n693), .ZN(n989) );
  INV_X1 U783 ( .A(KEYINPUT104), .ZN(n703) );
  INV_X1 U784 ( .A(n694), .ZN(n696) );
  NAND2_X1 U785 ( .A1(n696), .A2(n695), .ZN(n738) );
  INV_X1 U786 ( .A(G2072), .ZN(n955) );
  NOR2_X1 U787 ( .A1(n738), .A2(n955), .ZN(n699) );
  XOR2_X1 U788 ( .A(KEYINPUT103), .B(KEYINPUT27), .Z(n697) );
  XNOR2_X1 U789 ( .A(KEYINPUT102), .B(n697), .ZN(n698) );
  XNOR2_X1 U790 ( .A(n699), .B(n698), .ZN(n701) );
  NAND2_X1 U791 ( .A1(n738), .A2(G1956), .ZN(n700) );
  NAND2_X1 U792 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U793 ( .A(n703), .B(n702), .ZN(n722) );
  NOR2_X1 U794 ( .A1(n975), .A2(n722), .ZN(n704) );
  XOR2_X1 U795 ( .A(n704), .B(KEYINPUT28), .Z(n726) );
  NAND2_X1 U796 ( .A1(G1348), .A2(n738), .ZN(n706) );
  INV_X1 U797 ( .A(n738), .ZN(n729) );
  NAND2_X1 U798 ( .A1(G2067), .A2(n729), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n718) );
  NAND2_X1 U800 ( .A1(n718), .A2(n849), .ZN(n717) );
  XOR2_X1 U801 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n708) );
  NAND2_X1 U802 ( .A1(G1996), .A2(n708), .ZN(n707) );
  OR2_X1 U803 ( .A1(n738), .A2(n707), .ZN(n711) );
  INV_X1 U804 ( .A(G1996), .ZN(n954) );
  NOR2_X1 U805 ( .A1(n738), .A2(n954), .ZN(n709) );
  OR2_X1 U806 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U807 ( .A1(n711), .A2(n710), .ZN(n714) );
  AND2_X1 U808 ( .A1(n738), .A2(G1341), .ZN(n712) );
  NOR2_X1 U809 ( .A1(n712), .A2(n979), .ZN(n713) );
  AND2_X1 U810 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U811 ( .A(n715), .B(KEYINPUT65), .Z(n716) );
  NAND2_X1 U812 ( .A1(n717), .A2(n716), .ZN(n720) );
  OR2_X1 U813 ( .A1(n718), .A2(n849), .ZN(n719) );
  NAND2_X1 U814 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U815 ( .A(n721), .B(KEYINPUT105), .ZN(n724) );
  NAND2_X1 U816 ( .A1(n975), .A2(n722), .ZN(n723) );
  NAND2_X1 U817 ( .A1(n724), .A2(n723), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n726), .A2(n725), .ZN(n728) );
  XNOR2_X1 U819 ( .A(n728), .B(n727), .ZN(n735) );
  XOR2_X1 U820 ( .A(G2078), .B(KEYINPUT25), .Z(n960) );
  NOR2_X1 U821 ( .A1(n960), .A2(n738), .ZN(n731) );
  NOR2_X1 U822 ( .A1(n729), .A2(G1961), .ZN(n730) );
  NOR2_X1 U823 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U824 ( .A(KEYINPUT100), .B(n732), .ZN(n736) );
  NOR2_X1 U825 ( .A1(G301), .A2(n736), .ZN(n733) );
  XNOR2_X1 U826 ( .A(n733), .B(KEYINPUT101), .ZN(n734) );
  NAND2_X1 U827 ( .A1(n735), .A2(n734), .ZN(n747) );
  AND2_X1 U828 ( .A1(G301), .A2(n736), .ZN(n737) );
  XNOR2_X1 U829 ( .A(n737), .B(KEYINPUT106), .ZN(n744) );
  NAND2_X1 U830 ( .A1(n738), .A2(G8), .ZN(n739) );
  XNOR2_X1 U831 ( .A(n739), .B(KEYINPUT96), .ZN(n769) );
  NOR2_X1 U832 ( .A1(n769), .A2(G1966), .ZN(n760) );
  NOR2_X1 U833 ( .A1(G2084), .A2(n738), .ZN(n755) );
  NOR2_X1 U834 ( .A1(n760), .A2(n755), .ZN(n740) );
  NAND2_X1 U835 ( .A1(G8), .A2(n740), .ZN(n741) );
  XNOR2_X1 U836 ( .A(KEYINPUT30), .B(n741), .ZN(n742) );
  NOR2_X1 U837 ( .A1(n742), .A2(G168), .ZN(n743) );
  NOR2_X1 U838 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U839 ( .A(KEYINPUT31), .B(n745), .Z(n746) );
  NAND2_X1 U840 ( .A1(n757), .A2(G286), .ZN(n752) );
  NOR2_X1 U841 ( .A1(n769), .A2(G1971), .ZN(n749) );
  NOR2_X1 U842 ( .A1(G2090), .A2(n738), .ZN(n748) );
  NOR2_X1 U843 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U844 ( .A1(n750), .A2(G303), .ZN(n751) );
  NAND2_X1 U845 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U846 ( .A1(G8), .A2(n753), .ZN(n754) );
  XOR2_X1 U847 ( .A(KEYINPUT32), .B(n754), .Z(n763) );
  NAND2_X1 U848 ( .A1(G8), .A2(n755), .ZN(n756) );
  XOR2_X1 U849 ( .A(KEYINPUT99), .B(n756), .Z(n758) );
  NAND2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U851 ( .A(KEYINPUT107), .B(n761), .Z(n762) );
  NOR2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n782) );
  OR2_X1 U853 ( .A1(n989), .A2(n782), .ZN(n766) );
  NAND2_X1 U854 ( .A1(G1976), .A2(G288), .ZN(n982) );
  NOR2_X1 U855 ( .A1(n769), .A2(n764), .ZN(n765) );
  INV_X1 U856 ( .A(KEYINPUT33), .ZN(n767) );
  AND2_X1 U857 ( .A1(n768), .A2(KEYINPUT33), .ZN(n770) );
  INV_X1 U858 ( .A(n769), .ZN(n783) );
  NAND2_X1 U859 ( .A1(n770), .A2(n783), .ZN(n772) );
  XNOR2_X1 U860 ( .A(G1981), .B(G305), .ZN(n995) );
  NAND2_X1 U861 ( .A1(n773), .A2(n521), .ZN(n779) );
  NOR2_X1 U862 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U863 ( .A(KEYINPUT24), .B(KEYINPUT98), .Z(n774) );
  XNOR2_X1 U864 ( .A(KEYINPUT97), .B(n774), .ZN(n775) );
  XNOR2_X1 U865 ( .A(n776), .B(n775), .ZN(n777) );
  NAND2_X1 U866 ( .A1(n777), .A2(n783), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n786) );
  NAND2_X1 U868 ( .A1(G8), .A2(G166), .ZN(n780) );
  NOR2_X1 U869 ( .A1(G2090), .A2(n780), .ZN(n781) );
  NOR2_X1 U870 ( .A1(n782), .A2(n781), .ZN(n784) );
  NOR2_X1 U871 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U873 ( .A1(n788), .A2(n787), .ZN(n826) );
  NAND2_X1 U874 ( .A1(n903), .A2(G117), .ZN(n789) );
  XNOR2_X1 U875 ( .A(KEYINPUT91), .B(n789), .ZN(n792) );
  NAND2_X1 U876 ( .A1(n902), .A2(G129), .ZN(n790) );
  XOR2_X1 U877 ( .A(KEYINPUT90), .B(n790), .Z(n791) );
  NOR2_X1 U878 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U879 ( .A(KEYINPUT92), .B(n793), .Z(n797) );
  NAND2_X1 U880 ( .A1(G105), .A2(n906), .ZN(n794) );
  XNOR2_X1 U881 ( .A(n794), .B(KEYINPUT38), .ZN(n795) );
  XNOR2_X1 U882 ( .A(KEYINPUT93), .B(n795), .ZN(n796) );
  NOR2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n799) );
  NAND2_X1 U884 ( .A1(G141), .A2(n613), .ZN(n798) );
  NAND2_X1 U885 ( .A1(n799), .A2(n798), .ZN(n912) );
  NAND2_X1 U886 ( .A1(G1996), .A2(n912), .ZN(n800) );
  XNOR2_X1 U887 ( .A(n800), .B(KEYINPUT94), .ZN(n809) );
  NAND2_X1 U888 ( .A1(n906), .A2(G95), .ZN(n802) );
  NAND2_X1 U889 ( .A1(G131), .A2(n613), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U891 ( .A(KEYINPUT89), .B(n803), .ZN(n807) );
  NAND2_X1 U892 ( .A1(G119), .A2(n902), .ZN(n805) );
  NAND2_X1 U893 ( .A1(G107), .A2(n903), .ZN(n804) );
  AND2_X1 U894 ( .A1(n805), .A2(n804), .ZN(n806) );
  NAND2_X1 U895 ( .A1(n807), .A2(n806), .ZN(n898) );
  NAND2_X1 U896 ( .A1(G1991), .A2(n898), .ZN(n808) );
  NAND2_X1 U897 ( .A1(n809), .A2(n808), .ZN(n930) );
  NAND2_X1 U898 ( .A1(n930), .A2(n834), .ZN(n810) );
  XNOR2_X1 U899 ( .A(n810), .B(KEYINPUT95), .ZN(n830) );
  INV_X1 U900 ( .A(n830), .ZN(n824) );
  NAND2_X1 U901 ( .A1(G128), .A2(n902), .ZN(n812) );
  NAND2_X1 U902 ( .A1(G116), .A2(n903), .ZN(n811) );
  NAND2_X1 U903 ( .A1(n812), .A2(n811), .ZN(n813) );
  XNOR2_X1 U904 ( .A(n813), .B(KEYINPUT35), .ZN(n818) );
  NAND2_X1 U905 ( .A1(n906), .A2(G104), .ZN(n815) );
  NAND2_X1 U906 ( .A1(G140), .A2(n613), .ZN(n814) );
  NAND2_X1 U907 ( .A1(n815), .A2(n814), .ZN(n816) );
  XOR2_X1 U908 ( .A(KEYINPUT34), .B(n816), .Z(n817) );
  NAND2_X1 U909 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U910 ( .A(n819), .B(KEYINPUT36), .ZN(n899) );
  XOR2_X1 U911 ( .A(KEYINPUT37), .B(G2067), .Z(n820) );
  NOR2_X1 U912 ( .A1(n899), .A2(n820), .ZN(n932) );
  NAND2_X1 U913 ( .A1(n834), .A2(n932), .ZN(n836) );
  INV_X1 U914 ( .A(n836), .ZN(n823) );
  NAND2_X1 U915 ( .A1(n899), .A2(n820), .ZN(n821) );
  XOR2_X1 U916 ( .A(KEYINPUT88), .B(n821), .Z(n946) );
  NAND2_X1 U917 ( .A1(n946), .A2(n834), .ZN(n822) );
  OR2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n827) );
  AND2_X1 U919 ( .A1(n824), .A2(n827), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n841) );
  INV_X1 U921 ( .A(n827), .ZN(n839) );
  NOR2_X1 U922 ( .A1(G1996), .A2(n912), .ZN(n927) );
  NOR2_X1 U923 ( .A1(G1986), .A2(G290), .ZN(n828) );
  NOR2_X1 U924 ( .A1(G1991), .A2(n898), .ZN(n934) );
  NOR2_X1 U925 ( .A1(n828), .A2(n934), .ZN(n829) );
  NOR2_X1 U926 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U927 ( .A1(n927), .A2(n831), .ZN(n832) );
  XNOR2_X1 U928 ( .A(n832), .B(KEYINPUT39), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n833), .B(KEYINPUT108), .ZN(n835) );
  NAND2_X1 U930 ( .A1(n835), .A2(n834), .ZN(n837) );
  AND2_X1 U931 ( .A1(n837), .A2(n836), .ZN(n838) );
  OR2_X1 U932 ( .A1(n839), .A2(n838), .ZN(n840) );
  NAND2_X1 U933 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U934 ( .A(n842), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U935 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U936 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U937 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U938 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U939 ( .A1(n846), .A2(n845), .ZN(G188) );
  INV_X1 U941 ( .A(G132), .ZN(G219) );
  INV_X1 U942 ( .A(G120), .ZN(G236) );
  INV_X1 U943 ( .A(G82), .ZN(G220) );
  INV_X1 U944 ( .A(G69), .ZN(G235) );
  NOR2_X1 U945 ( .A1(n848), .A2(n847), .ZN(G325) );
  INV_X1 U946 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U947 ( .A(n979), .B(KEYINPUT116), .ZN(n851) );
  XNOR2_X1 U948 ( .A(G171), .B(n849), .ZN(n850) );
  XNOR2_X1 U949 ( .A(n851), .B(n850), .ZN(n854) );
  XOR2_X1 U950 ( .A(G286), .B(n852), .Z(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(n855) );
  NOR2_X1 U952 ( .A1(G37), .A2(n855), .ZN(G397) );
  XOR2_X1 U953 ( .A(G2678), .B(KEYINPUT43), .Z(n857) );
  XNOR2_X1 U954 ( .A(KEYINPUT42), .B(KEYINPUT109), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U956 ( .A(KEYINPUT110), .B(G2072), .Z(n859) );
  XNOR2_X1 U957 ( .A(G2067), .B(G2090), .ZN(n858) );
  XNOR2_X1 U958 ( .A(n859), .B(n858), .ZN(n860) );
  XOR2_X1 U959 ( .A(n861), .B(n860), .Z(n863) );
  XNOR2_X1 U960 ( .A(G2096), .B(G2100), .ZN(n862) );
  XNOR2_X1 U961 ( .A(n863), .B(n862), .ZN(n865) );
  XOR2_X1 U962 ( .A(G2078), .B(G2084), .Z(n864) );
  XNOR2_X1 U963 ( .A(n865), .B(n864), .ZN(G227) );
  XOR2_X1 U964 ( .A(G1976), .B(G1956), .Z(n867) );
  XNOR2_X1 U965 ( .A(G1981), .B(G1966), .ZN(n866) );
  XNOR2_X1 U966 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U967 ( .A(G1991), .B(G1971), .Z(n869) );
  XNOR2_X1 U968 ( .A(G1961), .B(G1996), .ZN(n868) );
  XNOR2_X1 U969 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U970 ( .A(n871), .B(n870), .Z(n873) );
  XNOR2_X1 U971 ( .A(G2474), .B(KEYINPUT41), .ZN(n872) );
  XNOR2_X1 U972 ( .A(n873), .B(n872), .ZN(n875) );
  XOR2_X1 U973 ( .A(G1986), .B(KEYINPUT111), .Z(n874) );
  XNOR2_X1 U974 ( .A(n875), .B(n874), .ZN(G229) );
  NAND2_X1 U975 ( .A1(G124), .A2(n902), .ZN(n876) );
  XNOR2_X1 U976 ( .A(n876), .B(KEYINPUT44), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n877), .B(KEYINPUT112), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G112), .A2(n903), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n883) );
  NAND2_X1 U980 ( .A1(n906), .A2(G100), .ZN(n881) );
  NAND2_X1 U981 ( .A1(G136), .A2(n613), .ZN(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  NOR2_X1 U983 ( .A1(n883), .A2(n882), .ZN(G162) );
  NAND2_X1 U984 ( .A1(n902), .A2(G127), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n884), .B(KEYINPUT114), .ZN(n886) );
  NAND2_X1 U986 ( .A1(G115), .A2(n903), .ZN(n885) );
  NAND2_X1 U987 ( .A1(n886), .A2(n885), .ZN(n887) );
  XNOR2_X1 U988 ( .A(n887), .B(KEYINPUT47), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G103), .A2(n906), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n892) );
  NAND2_X1 U991 ( .A1(G139), .A2(n613), .ZN(n890) );
  XNOR2_X1 U992 ( .A(KEYINPUT113), .B(n890), .ZN(n891) );
  NOR2_X1 U993 ( .A1(n892), .A2(n891), .ZN(n893) );
  XOR2_X1 U994 ( .A(KEYINPUT115), .B(n893), .Z(n937) );
  XOR2_X1 U995 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n895) );
  XNOR2_X1 U996 ( .A(G162), .B(n933), .ZN(n894) );
  XNOR2_X1 U997 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U998 ( .A(n937), .B(n896), .Z(n897) );
  XNOR2_X1 U999 ( .A(n898), .B(n897), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n899), .B(G160), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n916) );
  NAND2_X1 U1002 ( .A1(G130), .A2(n902), .ZN(n905) );
  NAND2_X1 U1003 ( .A1(G118), .A2(n903), .ZN(n904) );
  NAND2_X1 U1004 ( .A1(n905), .A2(n904), .ZN(n911) );
  NAND2_X1 U1005 ( .A1(n906), .A2(G106), .ZN(n908) );
  NAND2_X1 U1006 ( .A1(G142), .A2(n613), .ZN(n907) );
  NAND2_X1 U1007 ( .A1(n908), .A2(n907), .ZN(n909) );
  XOR2_X1 U1008 ( .A(n909), .B(KEYINPUT45), .Z(n910) );
  NOR2_X1 U1009 ( .A1(n911), .A2(n910), .ZN(n913) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1011 ( .A(G164), .B(n914), .Z(n915) );
  XNOR2_X1 U1012 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n917), .ZN(G395) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n925), .ZN(n922) );
  NOR2_X1 U1015 ( .A1(G227), .A2(G229), .ZN(n918) );
  XOR2_X1 U1016 ( .A(KEYINPUT49), .B(n918), .Z(n919) );
  XNOR2_X1 U1017 ( .A(n919), .B(KEYINPUT117), .ZN(n920) );
  NOR2_X1 U1018 ( .A1(G397), .A2(n920), .ZN(n921) );
  NAND2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  NOR2_X1 U1020 ( .A1(n923), .A2(G395), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(n924), .B(KEYINPUT118), .ZN(G308) );
  INV_X1 U1022 ( .A(G308), .ZN(G225) );
  INV_X1 U1023 ( .A(n925), .ZN(G319) );
  INV_X1 U1024 ( .A(G96), .ZN(G221) );
  INV_X1 U1025 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1026 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n1034) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n926) );
  NOR2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n928) );
  XNOR2_X1 U1029 ( .A(n928), .B(KEYINPUT51), .ZN(n929) );
  NOR2_X1 U1030 ( .A1(n930), .A2(n929), .ZN(n944) );
  XOR2_X1 U1031 ( .A(G2084), .B(G160), .Z(n931) );
  NOR2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n942) );
  XOR2_X1 U1035 ( .A(G164), .B(G2078), .Z(n939) );
  XNOR2_X1 U1036 ( .A(n955), .B(n937), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1038 ( .A(KEYINPUT50), .B(n940), .Z(n941) );
  NOR2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(n944), .A2(n943), .ZN(n945) );
  NOR2_X1 U1041 ( .A1(n946), .A2(n945), .ZN(n947) );
  XOR2_X1 U1042 ( .A(KEYINPUT52), .B(n947), .Z(n948) );
  XNOR2_X1 U1043 ( .A(KEYINPUT119), .B(n948), .ZN(n950) );
  INV_X1 U1044 ( .A(KEYINPUT55), .ZN(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1046 ( .A1(n951), .A2(G29), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(KEYINPUT120), .B(n952), .ZN(n1032) );
  XOR2_X1 U1048 ( .A(G2067), .B(G26), .Z(n953) );
  NAND2_X1 U1049 ( .A1(n953), .A2(G28), .ZN(n959) );
  XNOR2_X1 U1050 ( .A(n954), .B(G32), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n955), .B(G33), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n964) );
  XNOR2_X1 U1054 ( .A(n960), .B(G27), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(G1991), .B(G25), .ZN(n961) );
  NOR2_X1 U1056 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1057 ( .A1(n964), .A2(n963), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(n965), .B(KEYINPUT53), .ZN(n968) );
  XOR2_X1 U1059 ( .A(G2084), .B(G34), .Z(n966) );
  XNOR2_X1 U1060 ( .A(KEYINPUT54), .B(n966), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(G35), .B(G2090), .ZN(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1064 ( .A(KEYINPUT55), .B(n971), .ZN(n973) );
  INV_X1 U1065 ( .A(G29), .ZN(n972) );
  NAND2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n974), .A2(G11), .ZN(n1030) );
  XNOR2_X1 U1068 ( .A(G16), .B(KEYINPUT56), .ZN(n1001) );
  XNOR2_X1 U1069 ( .A(n975), .B(G1956), .ZN(n976) );
  XNOR2_X1 U1070 ( .A(n976), .B(KEYINPUT122), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(G1971), .A2(G303), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n978), .A2(n977), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(G1341), .B(n979), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n983) );
  NAND2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n993) );
  XNOR2_X1 U1076 ( .A(G171), .B(G1961), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(n984), .B(G1348), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(KEYINPUT121), .B(n987), .ZN(n991) );
  NOR2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n998) );
  XOR2_X1 U1083 ( .A(G168), .B(G1966), .Z(n994) );
  NOR2_X1 U1084 ( .A1(n995), .A2(n994), .ZN(n996) );
  XOR2_X1 U1085 ( .A(KEYINPUT57), .B(n996), .Z(n997) );
  NAND2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  XOR2_X1 U1087 ( .A(KEYINPUT123), .B(n999), .Z(n1000) );
  NAND2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1028) );
  INV_X1 U1089 ( .A(G16), .ZN(n1026) );
  XNOR2_X1 U1090 ( .A(G1348), .B(KEYINPUT59), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(n1002), .B(G4), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(G1956), .B(G20), .ZN(n1004) );
  XNOR2_X1 U1093 ( .A(G19), .B(G1341), .ZN(n1003) );
  NOR2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1009) );
  XOR2_X1 U1096 ( .A(KEYINPUT125), .B(G1981), .Z(n1007) );
  XNOR2_X1 U1097 ( .A(G6), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1099 ( .A(KEYINPUT60), .B(n1010), .Z(n1012) );
  XNOR2_X1 U1100 ( .A(G1966), .B(G21), .ZN(n1011) );
  NOR2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(n1013), .B(KEYINPUT126), .ZN(n1016) );
  XOR2_X1 U1103 ( .A(G1961), .B(G5), .Z(n1014) );
  XNOR2_X1 U1104 ( .A(KEYINPUT124), .B(n1014), .ZN(n1015) );
  NAND2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1023) );
  XNOR2_X1 U1106 ( .A(G1971), .B(G22), .ZN(n1018) );
  XNOR2_X1 U1107 ( .A(G23), .B(G1976), .ZN(n1017) );
  NOR2_X1 U1108 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  XOR2_X1 U1109 ( .A(G1986), .B(G24), .Z(n1019) );
  NAND2_X1 U1110 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1111 ( .A(KEYINPUT58), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1112 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1114 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1115 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NOR2_X1 U1116 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NAND2_X1 U1117 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  XNOR2_X1 U1118 ( .A(n1034), .B(n1033), .ZN(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

