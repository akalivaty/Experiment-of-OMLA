//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n768, new_n769, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n848, new_n849, new_n850,
    new_n851, new_n852, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956, new_n957;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n203));
  XNOR2_X1  g002(.A(G211gat), .B(G218gat), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  XNOR2_X1  g005(.A(KEYINPUT71), .B(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G197gat), .B(G204gat), .ZN(new_n210));
  AOI211_X1 g009(.A(new_n203), .B(new_n205), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G211gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT71), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT71), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G211gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n208), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n210), .B1(new_n216), .B2(KEYINPUT22), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n204), .B1(new_n217), .B2(KEYINPUT72), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n211), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT3), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  INV_X1    g020(.A(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT2), .ZN(new_n224));
  NAND2_X1  g023(.A1(G141gat), .A2(G148gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(G162gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G155gat), .ZN(new_n228));
  INV_X1    g027(.A(G155gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n229), .A2(G162gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n229), .A2(KEYINPUT76), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT76), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G155gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n224), .B1(new_n236), .B2(G162gat), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n223), .A2(new_n228), .A3(new_n230), .A4(new_n225), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n220), .B(new_n232), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT77), .ZN(new_n240));
  XNOR2_X1  g039(.A(KEYINPUT76), .B(G155gat), .ZN(new_n241));
  OAI21_X1  g040(.A(KEYINPUT2), .B1(new_n241), .B2(new_n227), .ZN(new_n242));
  INV_X1    g041(.A(new_n238), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT77), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n244), .A2(new_n245), .A3(new_n220), .A4(new_n232), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n240), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n219), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n242), .A2(new_n243), .B1(new_n226), .B2(new_n231), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n217), .A2(new_n205), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n209), .A2(new_n210), .A3(new_n204), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n248), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n250), .B1(new_n254), .B2(new_n220), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n202), .B1(new_n249), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G22gat), .ZN(new_n257));
  XOR2_X1   g056(.A(G197gat), .B(G204gat), .Z(new_n258));
  NOR2_X1   g057(.A1(new_n214), .A2(G211gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n212), .A2(KEYINPUT71), .ZN(new_n260));
  OAI21_X1  g059(.A(G218gat), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n258), .B1(new_n261), .B2(new_n206), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n205), .B1(new_n262), .B2(new_n203), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT29), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n217), .A2(KEYINPUT72), .A3(new_n204), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT80), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT3), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n263), .A2(KEYINPUT80), .A3(new_n264), .A4(new_n265), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n250), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n248), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n271), .B1(new_n240), .B2(new_n246), .ZN(new_n272));
  OAI211_X1 g071(.A(G228gat), .B(G233gat), .C1(new_n272), .C2(new_n219), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n256), .B(new_n257), .C1(new_n270), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(KEYINPUT81), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n266), .A2(new_n267), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(new_n220), .A3(new_n269), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n232), .B1(new_n237), .B2(new_n238), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n249), .A2(new_n202), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT81), .ZN(new_n282));
  NAND4_X1  g081(.A1(new_n281), .A2(new_n282), .A3(new_n257), .A4(new_n256), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n284));
  INV_X1    g083(.A(new_n256), .ZN(new_n285));
  OAI21_X1  g084(.A(G22gat), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n275), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G78gat), .B(G106gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(KEYINPUT31), .B(G50gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(new_n288), .B(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(new_n290), .B(KEYINPUT79), .Z(new_n291));
  AND2_X1   g090(.A1(new_n274), .A2(new_n290), .ZN(new_n292));
  AOI22_X1  g091(.A1(new_n287), .A2(new_n291), .B1(new_n286), .B2(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n294));
  INV_X1    g093(.A(G120gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(G113gat), .ZN(new_n296));
  INV_X1    g095(.A(G113gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G120gat), .ZN(new_n298));
  AOI21_X1  g097(.A(KEYINPUT1), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G127gat), .B(G134gat), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n294), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G134gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(G127gat), .ZN(new_n303));
  INV_X1    g102(.A(G127gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G134gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(G113gat), .B(G120gat), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n306), .B(KEYINPUT68), .C1(new_n307), .C2(KEYINPUT1), .ZN(new_n308));
  OR3_X1    g107(.A1(new_n295), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT69), .B1(new_n295), .B2(G113gat), .ZN(new_n310));
  INV_X1    g109(.A(new_n298), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n306), .A2(KEYINPUT1), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n301), .A2(new_n308), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT4), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n314), .A2(KEYINPUT78), .A3(new_n315), .A4(new_n250), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT78), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n308), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n312), .A2(new_n313), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n250), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n317), .B1(new_n320), .B2(KEYINPUT4), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n314), .A2(new_n315), .A3(new_n250), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n316), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT5), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n314), .B1(KEYINPUT3), .B2(new_n278), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(new_n247), .ZN(new_n327));
  NAND2_X1  g126(.A1(G225gat), .A2(G233gat), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n324), .A2(new_n325), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n320), .A2(KEYINPUT4), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n322), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(new_n327), .A3(new_n328), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n318), .A2(new_n319), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n278), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n320), .ZN(new_n335));
  INV_X1    g134(.A(new_n328), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n325), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n329), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G1gat), .B(G29gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT0), .ZN(new_n341));
  XNOR2_X1  g140(.A(G57gat), .B(G85gat), .ZN(new_n342));
  XOR2_X1   g141(.A(new_n341), .B(new_n342), .Z(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT6), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n329), .A2(new_n338), .A3(new_n343), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n339), .A2(KEYINPUT6), .A3(new_n344), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n219), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT67), .ZN(new_n352));
  AND2_X1   g151(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(G176gat), .ZN(new_n356));
  AND2_X1   g155(.A1(new_n356), .A2(KEYINPUT23), .ZN(new_n357));
  INV_X1    g156(.A(G169gat), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(new_n356), .ZN(new_n359));
  NAND2_X1  g158(.A1(G169gat), .A2(G176gat), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT23), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n355), .A2(new_n357), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n363));
  OAI21_X1  g162(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(G183gat), .A2(G190gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n363), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT25), .B1(new_n362), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n361), .A2(new_n359), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT25), .ZN(new_n371));
  NOR2_X1   g170(.A1(G169gat), .A2(G176gat), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n371), .B1(new_n372), .B2(KEYINPUT23), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n370), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT66), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n363), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(G183gat), .ZN(new_n377));
  INV_X1    g176(.A(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g178(.A1(KEYINPUT66), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n376), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n366), .A2(KEYINPUT65), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT65), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n383), .A2(G183gat), .A3(G190gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT24), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n374), .B1(new_n381), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n352), .B1(new_n369), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT64), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n358), .ZN(new_n391));
  NAND2_X1  g190(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n391), .A2(KEYINPUT23), .A3(new_n356), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n370), .ZN(new_n394));
  INV_X1    g193(.A(new_n363), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n395), .B1(new_n366), .B2(new_n364), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n371), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n376), .A2(new_n379), .A3(new_n380), .ZN(new_n398));
  AOI21_X1  g197(.A(KEYINPUT24), .B1(new_n382), .B2(new_n384), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n370), .B(new_n373), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(new_n400), .A3(KEYINPUT67), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n377), .A2(KEYINPUT27), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT27), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(G183gat), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n402), .A2(new_n404), .A3(new_n378), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT28), .ZN(new_n406));
  XNOR2_X1  g205(.A(new_n405), .B(new_n406), .ZN(new_n407));
  OR2_X1    g206(.A1(new_n359), .A2(KEYINPUT26), .ZN(new_n408));
  INV_X1    g207(.A(new_n360), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n359), .B1(new_n409), .B2(KEYINPUT26), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n367), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n407), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G226gat), .A2(G233gat), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n389), .A2(new_n401), .A3(new_n412), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n397), .A2(new_n400), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n412), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n414), .A2(KEYINPUT29), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n351), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n389), .A2(new_n401), .A3(new_n412), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n271), .A2(new_n414), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n416), .A2(new_n412), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n421), .A2(new_n422), .B1(new_n423), .B2(new_n414), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n420), .B1(new_n351), .B2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT74), .ZN(new_n426));
  XNOR2_X1  g225(.A(G8gat), .B(G36gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(G64gat), .B(G92gat), .ZN(new_n428));
  XNOR2_X1  g227(.A(new_n427), .B(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n425), .A2(new_n426), .A3(KEYINPUT30), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n419), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n432), .A2(new_n219), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n401), .A2(new_n412), .ZN(new_n434));
  AOI21_X1  g233(.A(KEYINPUT67), .B1(new_n397), .B2(new_n400), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n422), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n423), .A2(new_n414), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(new_n351), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n433), .A2(new_n438), .A3(KEYINPUT30), .A4(new_n430), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT74), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n431), .A2(new_n440), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n425), .A2(new_n430), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n433), .A2(new_n438), .A3(new_n430), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT30), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT75), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n443), .A2(KEYINPUT75), .A3(new_n444), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n441), .B(new_n442), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n293), .B1(new_n350), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n314), .B1(new_n434), .B2(new_n435), .ZN(new_n449));
  AND2_X1   g248(.A1(G227gat), .A2(G233gat), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n389), .A2(new_n401), .A3(new_n412), .A4(new_n333), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT33), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(KEYINPUT32), .ZN(new_n455));
  XOR2_X1   g254(.A(G15gat), .B(G43gat), .Z(new_n456));
  XNOR2_X1  g255(.A(G71gat), .B(G99gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n454), .A2(new_n455), .A3(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n458), .ZN(new_n460));
  OAI211_X1 g259(.A(new_n452), .B(KEYINPUT32), .C1(new_n453), .C2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n450), .B1(new_n449), .B2(new_n451), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT34), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n464), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n462), .A2(new_n467), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n459), .A2(new_n465), .A3(new_n466), .A4(new_n461), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT70), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT36), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n462), .A2(new_n467), .ZN(new_n473));
  AOI22_X1  g272(.A1(new_n459), .A2(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT36), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  AND3_X1   g276(.A1(new_n448), .A2(new_n472), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n432), .A2(new_n351), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n436), .A2(new_n437), .A3(new_n219), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT82), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .A4(KEYINPUT37), .ZN(new_n482));
  XNOR2_X1  g281(.A(KEYINPUT83), .B(KEYINPUT37), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n433), .A2(new_n438), .A3(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n482), .A2(new_n429), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n479), .A2(new_n480), .A3(KEYINPUT37), .ZN(new_n486));
  AOI21_X1  g285(.A(KEYINPUT38), .B1(new_n486), .B2(KEYINPUT82), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT37), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n429), .B(new_n484), .C1(new_n425), .C2(new_n488), .ZN(new_n489));
  AOI22_X1  g288(.A1(new_n485), .A2(new_n487), .B1(new_n489), .B2(KEYINPUT38), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n490), .A2(new_n443), .A3(new_n349), .A4(new_n348), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n335), .A2(new_n336), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT39), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n315), .B1(new_n314), .B2(new_n250), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n322), .B1(new_n495), .B2(new_n317), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n496), .A2(new_n316), .B1(new_n247), .B2(new_n326), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n494), .B1(new_n497), .B2(new_n328), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n324), .A2(new_n327), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(new_n493), .A3(new_n336), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n498), .A2(new_n500), .A3(KEYINPUT40), .A4(new_n343), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n501), .A2(new_n345), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(new_n500), .A3(new_n343), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT40), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n442), .B1(new_n446), .B2(new_n445), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n431), .A2(new_n440), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n502), .B(new_n505), .C1(new_n506), .C2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n287), .A2(new_n291), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n292), .A2(new_n286), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n491), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n506), .A2(new_n507), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n348), .A2(new_n349), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n473), .A2(new_n474), .ZN(new_n515));
  NAND4_X1  g314(.A1(new_n511), .A2(new_n513), .A3(new_n514), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(KEYINPUT35), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n293), .A2(new_n470), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT35), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n518), .A2(new_n519), .A3(new_n513), .A4(new_n514), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n478), .A2(new_n512), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT14), .ZN(new_n522));
  INV_X1    g321(.A(G29gat), .ZN(new_n523));
  INV_X1    g322(.A(G36gat), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(KEYINPUT84), .ZN(new_n526));
  OAI21_X1  g325(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT84), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n526), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n530), .B1(G29gat), .B2(G36gat), .ZN(new_n531));
  XOR2_X1   g330(.A(G43gat), .B(G50gat), .Z(new_n532));
  INV_X1    g331(.A(KEYINPUT15), .ZN(new_n533));
  OR2_X1    g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OR2_X1    g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g334(.A1(new_n532), .A2(new_n533), .B1(new_n525), .B2(new_n527), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n534), .B(new_n536), .C1(new_n523), .C2(new_n524), .ZN(new_n537));
  AND2_X1   g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G15gat), .B(G22gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT16), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n539), .B1(new_n540), .B2(G1gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT85), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n541), .B(new_n542), .C1(G1gat), .C2(new_n539), .ZN(new_n543));
  INV_X1    g342(.A(G8gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n538), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n535), .A2(new_n537), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT17), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n535), .A2(new_n549), .A3(new_n537), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n546), .B1(new_n551), .B2(new_n545), .ZN(new_n552));
  NAND2_X1  g351(.A1(G229gat), .A2(G233gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g353(.A1(KEYINPUT86), .A2(KEYINPUT18), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n552), .B(new_n553), .C1(KEYINPUT86), .C2(KEYINPUT18), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n546), .A2(KEYINPUT88), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT88), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n559), .B1(new_n538), .B2(new_n545), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n546), .B2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(KEYINPUT87), .B(KEYINPUT13), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n562), .B(new_n553), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n556), .A2(new_n557), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G113gat), .B(G141gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n566), .B(KEYINPUT11), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(new_n358), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(G197gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(KEYINPUT12), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n565), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n556), .A2(new_n557), .A3(new_n564), .A4(new_n570), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n521), .A2(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(G183gat), .B(G211gat), .Z(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT91), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(G71gat), .B(G78gat), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n581), .A2(KEYINPUT89), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n583));
  NOR2_X1   g382(.A1(G57gat), .A2(G64gat), .ZN(new_n584));
  AND2_X1   g383(.A1(G57gat), .A2(G64gat), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n581), .A2(KEYINPUT89), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT90), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(new_n586), .A2(new_n581), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT21), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G231gat), .ZN(new_n595));
  INV_X1    g394(.A(G233gat), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n592), .B(new_n593), .C1(new_n595), .C2(new_n596), .ZN(new_n599));
  XNOR2_X1  g398(.A(G127gat), .B(G155gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n600), .B1(new_n598), .B2(new_n599), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n580), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n605), .A2(new_n601), .A3(new_n579), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n545), .B1(new_n592), .B2(new_n593), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n607), .B1(new_n604), .B2(new_n606), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n577), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n610), .ZN(new_n612));
  INV_X1    g411(.A(new_n577), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G134gat), .B(G162gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n615), .B(KEYINPUT93), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G85gat), .A2(G92gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(new_n618), .B(KEYINPUT7), .ZN(new_n619));
  INV_X1    g418(.A(G99gat), .ZN(new_n620));
  INV_X1    g419(.A(G106gat), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT8), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n619), .B(new_n622), .C1(G85gat), .C2(G92gat), .ZN(new_n623));
  XOR2_X1   g422(.A(G99gat), .B(G106gat), .Z(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n551), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(G232gat), .A2(G233gat), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n628), .A2(KEYINPUT41), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n629), .B1(new_n547), .B2(new_n625), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT94), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI211_X1 g431(.A(KEYINPUT94), .B(new_n629), .C1(new_n547), .C2(new_n625), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n627), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G190gat), .B(G218gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n635), .ZN(new_n637));
  OAI211_X1 g436(.A(new_n627), .B(new_n637), .C1(new_n632), .C2(new_n633), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n628), .A2(KEYINPUT41), .ZN(new_n639));
  XNOR2_X1  g438(.A(new_n639), .B(KEYINPUT92), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n636), .A2(new_n638), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n641), .B1(new_n636), .B2(new_n638), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n617), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n636), .A2(new_n638), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n640), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n636), .A2(new_n638), .A3(new_n641), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n646), .A2(new_n616), .A3(new_n647), .ZN(new_n648));
  AOI22_X1  g447(.A1(new_n611), .A2(new_n614), .B1(new_n644), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n592), .B(new_n626), .ZN(new_n650));
  NAND2_X1  g449(.A1(G230gat), .A2(G233gat), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT95), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n592), .A2(new_n626), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n625), .B1(new_n590), .B2(new_n591), .ZN(new_n656));
  OR3_X1    g455(.A1(new_n655), .A2(new_n656), .A3(KEYINPUT10), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(KEYINPUT10), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n652), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(KEYINPUT96), .B1(new_n654), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(G176gat), .B(G204gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n663), .ZN(new_n665));
  OAI211_X1 g464(.A(KEYINPUT96), .B(new_n665), .C1(new_n654), .C2(new_n659), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n649), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n576), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n514), .A2(KEYINPUT97), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n514), .A2(KEYINPUT97), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g474(.A1(new_n670), .A2(new_n447), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT98), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT16), .B1(new_n677), .B2(KEYINPUT42), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT42), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n540), .A2(new_n679), .A3(KEYINPUT98), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n676), .B1(new_n678), .B2(new_n680), .ZN(new_n681));
  OR2_X1    g480(.A1(new_n681), .A2(new_n544), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n544), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n676), .A2(new_n679), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n682), .A2(new_n683), .A3(new_n684), .ZN(G1325gat));
  NOR3_X1   g484(.A1(new_n669), .A2(G15gat), .A3(new_n470), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n477), .A2(new_n472), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n686), .B1(G15gat), .B2(new_n688), .ZN(new_n689));
  XOR2_X1   g488(.A(new_n689), .B(KEYINPUT99), .Z(G1326gat));
  NOR2_X1   g489(.A1(new_n669), .A2(new_n511), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  INV_X1    g492(.A(new_n667), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n614), .A2(new_n611), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n644), .A2(new_n648), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n694), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n576), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n698), .A2(new_n523), .A3(new_n673), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT100), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT45), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n695), .A2(KEYINPUT101), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT101), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n614), .A2(new_n611), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n705), .A2(new_n574), .A3(new_n667), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT102), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n517), .A2(new_n520), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n512), .A2(new_n472), .A3(new_n477), .A4(new_n448), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n696), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n707), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g511(.A(KEYINPUT102), .B(KEYINPUT44), .C1(new_n521), .C2(new_n696), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT103), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n521), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n708), .A2(new_n709), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(KEYINPUT103), .ZN(new_n718));
  AND2_X1   g517(.A1(new_n644), .A2(new_n648), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n716), .A2(new_n718), .A3(new_n711), .A4(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n706), .B1(new_n714), .B2(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n721), .A2(new_n673), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n701), .B1(new_n523), .B2(new_n722), .ZN(G1328gat));
  NAND3_X1  g522(.A1(new_n698), .A2(new_n524), .A3(new_n447), .ZN(new_n724));
  XOR2_X1   g523(.A(new_n724), .B(KEYINPUT46), .Z(new_n725));
  AND2_X1   g524(.A1(new_n721), .A2(new_n447), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n524), .B2(new_n726), .ZN(G1329gat));
  INV_X1    g526(.A(G43gat), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n698), .A2(new_n728), .A3(new_n515), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n721), .A2(new_n687), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n730), .B2(new_n728), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT47), .B1(new_n729), .B2(KEYINPUT104), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1330gat));
  INV_X1    g532(.A(G50gat), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n576), .A2(new_n734), .A3(new_n293), .A4(new_n697), .ZN(new_n735));
  AOI211_X1 g534(.A(new_n511), .B(new_n706), .C1(new_n714), .C2(new_n720), .ZN(new_n736));
  OAI211_X1 g535(.A(KEYINPUT48), .B(new_n735), .C1(new_n736), .C2(new_n734), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT106), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n735), .B(new_n738), .ZN(new_n739));
  AOI21_X1  g538(.A(new_n734), .B1(new_n721), .B2(new_n293), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n739), .B1(new_n740), .B2(KEYINPUT105), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT105), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n736), .B2(new_n734), .ZN(new_n743));
  AOI211_X1 g542(.A(KEYINPUT107), .B(KEYINPUT48), .C1(new_n741), .C2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n714), .A2(new_n720), .ZN(new_n746));
  INV_X1    g545(.A(new_n706), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n746), .A2(new_n293), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n748), .A2(KEYINPUT105), .A3(G50gat), .ZN(new_n749));
  INV_X1    g548(.A(new_n739), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n743), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT48), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n745), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n737), .B1(new_n744), .B2(new_n753), .ZN(G1331gat));
  AND2_X1   g553(.A1(new_n716), .A2(new_n718), .ZN(new_n755));
  INV_X1    g554(.A(new_n695), .ZN(new_n756));
  NOR4_X1   g555(.A1(new_n756), .A2(new_n719), .A3(new_n574), .A4(new_n667), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n673), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n760), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g560(.A(new_n513), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n763), .B(new_n764), .Z(G1333gat));
  NAND3_X1  g564(.A1(new_n759), .A2(G71gat), .A3(new_n687), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n758), .A2(new_n470), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(G71gat), .B2(new_n767), .ZN(new_n768));
  XNOR2_X1  g567(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n768), .B(new_n769), .ZN(G1334gat));
  NAND2_X1  g569(.A1(new_n759), .A2(new_n293), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g571(.A1(new_n714), .A2(new_n720), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n756), .A2(new_n575), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n694), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(G85gat), .A3(new_n673), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n775), .A2(new_n710), .A3(KEYINPUT51), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT51), .B1(new_n775), .B2(new_n710), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n694), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(new_n673), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n778), .B1(G85gat), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT109), .ZN(G1336gat));
  NAND3_X1  g584(.A1(new_n777), .A2(G92gat), .A3(new_n447), .ZN(new_n786));
  INV_X1    g585(.A(G92gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(new_n781), .B2(new_n513), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n789), .B(KEYINPUT52), .Z(G1337gat));
  AOI21_X1  g589(.A(new_n620), .B1(new_n477), .B2(new_n472), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n781), .A2(new_n470), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n777), .A2(new_n791), .B1(new_n792), .B2(new_n620), .ZN(G1338gat));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n773), .A2(new_n511), .A3(new_n776), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n794), .B1(new_n795), .B2(new_n621), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT53), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OR3_X1    g597(.A1(new_n781), .A2(G106gat), .A3(new_n511), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n799), .B1(new_n795), .B2(new_n621), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n798), .B(new_n800), .ZN(G1339gat));
  INV_X1    g600(.A(new_n659), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n657), .A2(new_n658), .A3(new_n652), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(KEYINPUT54), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g603(.A(KEYINPUT112), .B(KEYINPUT54), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n665), .B1(new_n659), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n804), .A2(KEYINPUT55), .A3(new_n806), .ZN(new_n810));
  OR3_X1    g609(.A1(new_n654), .A2(new_n663), .A3(new_n659), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n574), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n561), .A2(new_n563), .B1(new_n553), .B2(new_n552), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(new_n569), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n664), .A2(new_n573), .A3(new_n666), .A4(new_n814), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n719), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n573), .A2(new_n814), .ZN(new_n818));
  NOR3_X1   g617(.A1(new_n817), .A2(new_n696), .A3(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n705), .B1(new_n816), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n695), .A2(new_n696), .A3(new_n575), .A4(new_n667), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(KEYINPUT111), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT111), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n649), .A2(new_n823), .A3(new_n575), .A4(new_n667), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n782), .B1(new_n820), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n826), .A2(new_n513), .A3(new_n518), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n828), .A2(KEYINPUT113), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT113), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n297), .B(new_n574), .C1(new_n829), .C2(new_n831), .ZN(new_n832));
  OAI21_X1  g631(.A(G113gat), .B1(new_n827), .B2(new_n575), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(G1340gat));
  OAI211_X1 g633(.A(new_n295), .B(new_n694), .C1(new_n829), .C2(new_n831), .ZN(new_n835));
  OAI21_X1  g634(.A(G120gat), .B1(new_n827), .B2(new_n667), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n835), .A2(KEYINPUT114), .A3(new_n836), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1341gat));
  AOI21_X1  g640(.A(G127gat), .B1(new_n828), .B2(new_n695), .ZN(new_n842));
  INV_X1    g641(.A(new_n705), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(G127gat), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT115), .B1(new_n827), .B2(new_n844), .ZN(new_n845));
  OR3_X1    g644(.A1(new_n827), .A2(KEYINPUT115), .A3(new_n844), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n842), .B1(new_n845), .B2(new_n846), .ZN(G1342gat));
  NOR2_X1   g646(.A1(new_n696), .A2(new_n447), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n826), .A2(new_n518), .A3(new_n848), .ZN(new_n849));
  OR3_X1    g648(.A1(new_n849), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT56), .B1(new_n849), .B2(G134gat), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(G134gat), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(G1343gat));
  NOR2_X1   g652(.A1(new_n687), .A2(new_n511), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT117), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n826), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n574), .A2(new_n221), .ZN(new_n857));
  XOR2_X1   g656(.A(new_n857), .B(KEYINPUT118), .Z(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n513), .A3(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT119), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n782), .A2(new_n687), .A3(new_n447), .ZN(new_n861));
  XOR2_X1   g660(.A(new_n861), .B(KEYINPUT116), .Z(new_n862));
  AOI21_X1  g661(.A(new_n511), .B1(new_n820), .B2(new_n825), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(KEYINPUT57), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n293), .A2(KEYINPUT57), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n756), .B1(new_n816), .B2(new_n819), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n865), .B1(new_n866), .B2(new_n825), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n574), .B(new_n862), .C1(new_n864), .C2(new_n867), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n868), .A2(G141gat), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT58), .B1(new_n860), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT58), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n868), .A2(KEYINPUT120), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(G141gat), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n868), .A2(KEYINPUT120), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n871), .B(new_n859), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n870), .A2(new_n875), .ZN(G1344gat));
  NOR2_X1   g675(.A1(new_n864), .A2(new_n867), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n862), .A2(new_n694), .ZN(new_n878));
  NOR3_X1   g677(.A1(new_n877), .A2(KEYINPUT59), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n856), .A2(new_n513), .ZN(new_n880));
  OAI21_X1  g679(.A(KEYINPUT59), .B1(new_n880), .B2(new_n667), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n879), .B1(new_n222), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n863), .A2(KEYINPUT121), .A3(KEYINPUT57), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT121), .B1(new_n863), .B2(KEYINPUT57), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n817), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n886), .A2(new_n719), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT122), .B1(new_n817), .B2(new_n696), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n818), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n756), .B1(new_n890), .B2(new_n816), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n821), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT57), .B1(new_n892), .B2(new_n293), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n885), .A2(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n894), .A2(new_n878), .ZN(new_n895));
  NAND2_X1  g694(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n882), .B1(new_n895), .B2(new_n896), .ZN(G1345gat));
  INV_X1    g696(.A(new_n862), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n877), .A2(new_n705), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n695), .A2(new_n241), .ZN(new_n900));
  OAI22_X1  g699(.A1(new_n899), .A2(new_n241), .B1(new_n880), .B2(new_n900), .ZN(G1346gat));
  NAND3_X1  g700(.A1(new_n856), .A2(new_n227), .A3(new_n848), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n877), .A2(new_n696), .A3(new_n898), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(new_n903), .B2(new_n227), .ZN(G1347gat));
  NAND2_X1  g703(.A1(new_n820), .A2(new_n825), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n673), .A2(new_n513), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT123), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n907), .A2(new_n518), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(G169gat), .B1(new_n909), .B2(new_n575), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n905), .A2(new_n906), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n518), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n574), .A2(new_n355), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(G1348gat));
  INV_X1    g713(.A(new_n912), .ZN(new_n915));
  AOI21_X1  g714(.A(G176gat), .B1(new_n915), .B2(new_n694), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n916), .A2(new_n917), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n909), .A2(new_n356), .A3(new_n667), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(G1349gat));
  OAI21_X1  g720(.A(G183gat), .B1(new_n909), .B2(new_n705), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n695), .A2(new_n402), .A3(new_n404), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n912), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n925));
  XOR2_X1   g724(.A(new_n924), .B(new_n925), .Z(G1350gat));
  NAND3_X1  g725(.A1(new_n915), .A2(new_n378), .A3(new_n719), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n905), .A2(new_n908), .A3(new_n719), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT61), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n928), .A2(new_n929), .A3(G190gat), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n928), .B2(G190gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n927), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n932), .B(new_n933), .ZN(G1351gat));
  NAND2_X1  g733(.A1(new_n911), .A2(new_n854), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(G197gat), .B1(new_n936), .B2(new_n574), .ZN(new_n937));
  INV_X1    g736(.A(new_n907), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n938), .A2(new_n687), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n894), .A2(new_n940), .ZN(new_n941));
  AND2_X1   g740(.A1(new_n574), .A2(G197gat), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n937), .B1(new_n941), .B2(new_n942), .ZN(G1352gat));
  NOR3_X1   g742(.A1(new_n935), .A2(G204gat), .A3(new_n667), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT62), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n894), .A2(new_n667), .A3(new_n940), .ZN(new_n946));
  INV_X1    g745(.A(G204gat), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(G1353gat));
  NAND3_X1  g747(.A1(new_n936), .A2(new_n207), .A3(new_n695), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n695), .B(new_n939), .C1(new_n885), .C2(new_n893), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n950), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT63), .B1(new_n950), .B2(G211gat), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(G1354gat));
  OAI21_X1  g752(.A(new_n208), .B1(new_n935), .B2(new_n696), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n954), .B(new_n955), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n696), .A2(new_n208), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n956), .B1(new_n941), .B2(new_n957), .ZN(G1355gat));
endmodule


