//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 1 1 1 1 0 1 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n617, new_n618, new_n621, new_n622, new_n624, new_n625, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1195, new_n1196, new_n1197,
    new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT68), .ZN(G217));
  NOR4_X1   g027(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT69), .Z(new_n459));
  AOI21_X1  g034(.A(new_n459), .B1(new_n454), .B2(G2106), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(KEYINPUT70), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT70), .ZN(new_n468));
  NAND2_X1  g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n464), .A2(new_n470), .A3(G125), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n461), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(G2105), .B1(new_n467), .B2(new_n469), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n466), .A2(G2105), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n474), .A2(G137), .B1(G101), .B2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n473), .A2(new_n477), .ZN(G160));
  OAI21_X1  g053(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n480), .B1(G112), .B2(new_n461), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT71), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n461), .B1(new_n467), .B2(new_n469), .ZN(new_n483));
  AOI22_X1  g058(.A1(G124), .A2(new_n483), .B1(new_n474), .B2(G136), .ZN(new_n484));
  AND2_X1   g059(.A1(new_n482), .A2(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n462), .C2(new_n463), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT72), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT72), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n486), .A2(new_n493), .A3(new_n490), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(G138), .ZN(new_n497));
  NOR3_X1   g072(.A1(new_n497), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n464), .A2(new_n470), .A3(new_n498), .ZN(new_n499));
  AOI22_X1  g074(.A1(new_n492), .A2(new_n494), .B1(new_n496), .B2(new_n499), .ZN(G164));
  NAND2_X1  g075(.A1(G75), .A2(G543), .ZN(new_n501));
  AND3_X1   g076(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n502));
  AOI21_X1  g077(.A(KEYINPUT5), .B1(KEYINPUT73), .B2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G62), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n501), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n506), .A2(G651), .B1(G50), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT74), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n514), .B1(new_n504), .B2(new_n509), .ZN(new_n515));
  OAI221_X1 g090(.A(KEYINPUT74), .B1(new_n507), .B2(new_n508), .C1(new_n502), .C2(new_n503), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n512), .B1(new_n513), .B2(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND2_X1  g094(.A1(new_n511), .A2(G51), .ZN(new_n520));
  OAI211_X1 g095(.A(G63), .B(G651), .C1(new_n502), .C2(new_n503), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(KEYINPUT75), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT7), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(KEYINPUT75), .ZN(new_n525));
  AND3_X1   g100(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AOI21_X1  g101(.A(new_n524), .B1(new_n523), .B2(new_n525), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n520), .B(new_n521), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  AND3_X1   g103(.A1(new_n515), .A2(G89), .A3(new_n516), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(G168));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  INV_X1    g106(.A(G77), .ZN(new_n532));
  OAI22_X1  g107(.A1(new_n504), .A2(new_n531), .B1(new_n532), .B2(new_n510), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT76), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI221_X1 g110(.A(KEYINPUT76), .B1(new_n532), .B2(new_n510), .C1(new_n504), .C2(new_n531), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n535), .A2(G651), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n511), .A2(G52), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n515), .A2(new_n516), .A3(G90), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(G171));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n504), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n544), .A2(G651), .B1(G43), .B2(new_n511), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n515), .A2(new_n516), .A3(G81), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n550));
  XOR2_X1   g125(.A(new_n550), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  XNOR2_X1  g130(.A(KEYINPUT78), .B(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n555), .B1(new_n504), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G651), .ZN(new_n558));
  INV_X1    g133(.A(G91), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n511), .A2(G53), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n560), .A2(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n562), .B1(new_n511), .B2(G53), .ZN(new_n563));
  OAI221_X1 g138(.A(new_n558), .B1(new_n517), .B2(new_n559), .C1(new_n561), .C2(new_n563), .ZN(G299));
  INV_X1    g139(.A(KEYINPUT79), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n540), .A2(new_n565), .ZN(new_n566));
  AND2_X1   g141(.A1(new_n539), .A2(new_n538), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n567), .A2(KEYINPUT79), .A3(new_n537), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  INV_X1    g144(.A(new_n569), .ZN(G301));
  INV_X1    g145(.A(G168), .ZN(G286));
  INV_X1    g146(.A(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n504), .A2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(G651), .A2(new_n573), .B1(new_n511), .B2(G49), .ZN(new_n574));
  INV_X1    g149(.A(G87), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n517), .ZN(G288));
  OAI21_X1  g151(.A(G61), .B1(new_n502), .B2(new_n503), .ZN(new_n577));
  AND3_X1   g152(.A1(KEYINPUT80), .A2(G73), .A3(G543), .ZN(new_n578));
  AOI21_X1  g153(.A(KEYINPUT80), .B1(G73), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g156(.A1(new_n581), .A2(G651), .B1(new_n511), .B2(G48), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n515), .A2(new_n516), .A3(G86), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(G305));
  NAND2_X1  g159(.A1(new_n511), .A2(G47), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n517), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT82), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(G72), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G60), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n504), .B2(new_n591), .ZN(new_n592));
  AND3_X1   g167(.A1(new_n592), .A2(KEYINPUT81), .A3(G651), .ZN(new_n593));
  AOI21_X1  g168(.A(KEYINPUT81), .B1(new_n592), .B2(G651), .ZN(new_n594));
  NOR2_X1   g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT82), .ZN(new_n596));
  OAI211_X1 g171(.A(new_n596), .B(new_n585), .C1(new_n517), .C2(new_n586), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n589), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(G290));
  AND2_X1   g175(.A1(new_n515), .A2(new_n516), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n601), .A2(KEYINPUT10), .A3(G92), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT10), .ZN(new_n603));
  INV_X1    g178(.A(G92), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n517), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n602), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g181(.A1(G79), .A2(G543), .ZN(new_n607));
  INV_X1    g182(.A(G66), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n504), .B2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n609), .A2(G651), .B1(G54), .B2(new_n511), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n611), .A2(G868), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(new_n569), .B2(G868), .ZN(G284));
  XOR2_X1   g188(.A(G284), .B(KEYINPUT83), .Z(G321));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n615));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NOR2_X1   g191(.A1(G168), .A2(new_n616), .ZN(new_n617));
  AOI211_X1 g192(.A(new_n615), .B(new_n617), .C1(new_n616), .C2(G299), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n618), .B1(new_n615), .B2(new_n617), .ZN(G297));
  AOI21_X1  g194(.A(new_n618), .B1(new_n615), .B2(new_n617), .ZN(G280));
  INV_X1    g195(.A(new_n611), .ZN(new_n621));
  INV_X1    g196(.A(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G860), .ZN(G148));
  NAND2_X1  g198(.A1(new_n547), .A2(new_n616), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n611), .A2(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(new_n616), .ZN(G323));
  XNOR2_X1  g201(.A(G323), .B(KEYINPUT11), .ZN(G282));
  AND2_X1   g202(.A1(new_n464), .A2(new_n470), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(new_n475), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT13), .Z(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  AOI22_X1  g209(.A1(G123), .A2(new_n483), .B1(new_n474), .B2(G135), .ZN(new_n635));
  NOR3_X1   g210(.A1(new_n461), .A2(KEYINPUT85), .A3(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(KEYINPUT85), .B1(new_n461), .B2(G111), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n637), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n635), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n634), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(new_n641), .B(KEYINPUT86), .Z(G156));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2427), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2430), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT15), .B(G2435), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(new_n646), .B2(new_n645), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2451), .B(G2454), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT16), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n648), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2443), .B(G2446), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT87), .ZN(G401));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT17), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2084), .B(G2090), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  NOR3_X1   g237(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT88), .Z(new_n664));
  NAND2_X1  g239(.A1(new_n660), .A2(new_n662), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n665), .B(new_n661), .C1(new_n659), .C2(new_n662), .ZN(new_n666));
  INV_X1    g241(.A(new_n661), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n667), .A2(new_n659), .A3(new_n662), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n666), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2096), .B(G2100), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(G227));
  XOR2_X1   g248(.A(G1971), .B(G1976), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT19), .ZN(new_n675));
  XOR2_X1   g250(.A(G1956), .B(G2474), .Z(new_n676));
  XOR2_X1   g251(.A(G1961), .B(G1966), .Z(new_n677));
  AND2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n676), .A2(new_n677), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  MUX2_X1   g258(.A(new_n683), .B(new_n682), .S(new_n675), .Z(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1991), .B(G1996), .Z(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n686), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n685), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n688), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  AND3_X1   g269(.A1(new_n689), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n694), .B1(new_n689), .B2(new_n693), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(G229));
  INV_X1    g272(.A(G16), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G22), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G166), .B2(new_n698), .ZN(new_n700));
  INV_X1    g275(.A(G1971), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(G6), .A2(G16), .ZN(new_n703));
  INV_X1    g278(.A(G305), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n703), .B1(new_n704), .B2(G16), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT32), .B(G1981), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(G16), .A2(G23), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT92), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G288), .B2(new_n698), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT33), .B(G1976), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n702), .A2(new_n707), .A3(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT34), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n599), .A2(G16), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G16), .B2(G24), .ZN(new_n716));
  INV_X1    g291(.A(G1986), .ZN(new_n717));
  OR2_X1    g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G25), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT90), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n474), .A2(G131), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n483), .A2(G119), .ZN(new_n723));
  OR2_X1    g298(.A1(G95), .A2(G2105), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n724), .B(G2104), .C1(G107), .C2(new_n461), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n722), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n721), .B1(new_n726), .B2(G29), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT35), .B(G1991), .Z(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT91), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n727), .B(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(new_n716), .B2(new_n717), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n714), .A2(new_n718), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(KEYINPUT93), .A2(KEYINPUT36), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n719), .A2(G35), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT98), .Z(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G162), .B2(new_n719), .ZN(new_n738));
  XNOR2_X1  g313(.A(KEYINPUT99), .B(KEYINPUT29), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n740), .A2(G2090), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n698), .A2(G20), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT23), .Z(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G299), .B2(G16), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(G1956), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n741), .A2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT100), .Z(new_n747));
  AND2_X1   g322(.A1(new_n719), .A2(G32), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n474), .A2(G141), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT96), .Z(new_n750));
  AND2_X1   g325(.A1(new_n475), .A2(G105), .ZN(new_n751));
  NAND3_X1  g326(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT26), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n751), .B(new_n753), .C1(G129), .C2(new_n483), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n748), .B1(new_n755), .B2(G29), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT27), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n758), .A2(G1996), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n719), .A2(G26), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT28), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n474), .A2(G140), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n483), .A2(G128), .ZN(new_n764));
  OR2_X1    g339(.A1(G104), .A2(G2105), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n765), .B(G2104), .C1(G116), .C2(new_n461), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n762), .B1(new_n768), .B2(new_n719), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT95), .B(G2067), .Z(new_n770));
  AND2_X1   g345(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT31), .B(G11), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT97), .B(G28), .Z(new_n774));
  AOI21_X1  g349(.A(G29), .B1(new_n774), .B2(KEYINPUT30), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(KEYINPUT30), .B2(new_n774), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n773), .B(new_n776), .C1(new_n639), .C2(new_n719), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n771), .A2(new_n772), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n719), .A2(G33), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n628), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(new_n461), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n782));
  XOR2_X1   g357(.A(new_n782), .B(KEYINPUT25), .Z(new_n783));
  NAND2_X1  g358(.A1(new_n474), .A2(G139), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n779), .B1(new_n786), .B2(new_n719), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n760), .B(new_n778), .C1(G2072), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n719), .A2(G27), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G164), .B2(new_n719), .ZN(new_n790));
  INV_X1    g365(.A(G2078), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(G2084), .ZN(new_n793));
  NAND2_X1  g368(.A1(G160), .A2(G29), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT24), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n795), .A2(G34), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n719), .B1(new_n795), .B2(G34), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI221_X1 g373(.A(new_n792), .B1(new_n793), .B2(new_n798), .C1(new_n740), .C2(G2090), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n787), .A2(G2072), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n698), .A2(G21), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G168), .B2(new_n698), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(G1966), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(G1966), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n798), .A2(new_n793), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n800), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  NOR3_X1   g381(.A1(new_n788), .A2(new_n799), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n698), .A2(G19), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n548), .B2(new_n698), .ZN(new_n809));
  INV_X1    g384(.A(G1341), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n758), .A2(new_n759), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n811), .B1(new_n812), .B2(G1996), .ZN(new_n813));
  NOR2_X1   g388(.A1(G4), .A2(G16), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT94), .Z(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n621), .B2(G16), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G1348), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n698), .A2(G5), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G171), .B2(new_n698), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(G1961), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n813), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n747), .A2(new_n807), .A3(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n822), .A2(KEYINPUT101), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(KEYINPUT101), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n734), .A2(new_n735), .B1(new_n823), .B2(new_n824), .ZN(G311));
  NAND2_X1  g400(.A1(new_n734), .A2(new_n735), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n823), .A2(new_n824), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(G150));
  NOR2_X1   g403(.A1(new_n611), .A2(new_n622), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n547), .A2(KEYINPUT103), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT103), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n545), .A2(new_n833), .A3(new_n546), .ZN(new_n834));
  NAND2_X1  g409(.A1(G80), .A2(G543), .ZN(new_n835));
  INV_X1    g410(.A(G67), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n504), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(G651), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n511), .A2(G55), .ZN(new_n839));
  INV_X1    g414(.A(G93), .ZN(new_n840));
  OAI211_X1 g415(.A(new_n838), .B(new_n839), .C1(new_n517), .C2(new_n840), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n832), .A2(new_n834), .A3(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n841), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n843), .A2(new_n548), .A3(new_n833), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n831), .B(new_n845), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT39), .ZN(new_n847));
  AOI21_X1  g422(.A(G860), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n847), .B2(new_n846), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(KEYINPUT104), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n841), .A2(G860), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT37), .Z(new_n852));
  NAND2_X1  g427(.A1(new_n850), .A2(new_n852), .ZN(G145));
  AOI22_X1  g428(.A1(G130), .A2(new_n483), .B1(new_n474), .B2(G142), .ZN(new_n854));
  OAI21_X1  g429(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n855));
  INV_X1    g430(.A(G118), .ZN(new_n856));
  AOI22_X1  g431(.A1(new_n855), .A2(KEYINPUT105), .B1(new_n856), .B2(G2105), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(KEYINPUT105), .B2(new_n855), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT106), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(new_n630), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n630), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n755), .A2(new_n767), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n755), .A2(new_n767), .ZN(new_n866));
  INV_X1    g441(.A(new_n726), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n755), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n869), .A2(new_n768), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n726), .B1(new_n870), .B2(new_n864), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n863), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n867), .B1(new_n865), .B2(new_n866), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n870), .A2(new_n726), .A3(new_n864), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n873), .A2(new_n862), .A3(new_n861), .A4(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n499), .A2(new_n496), .ZN(new_n876));
  INV_X1    g451(.A(new_n491), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n872), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n878), .B1(new_n872), .B2(new_n875), .ZN(new_n881));
  OAI22_X1  g456(.A1(new_n880), .A2(new_n881), .B1(new_n781), .B2(new_n785), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(new_n786), .A3(new_n879), .ZN(new_n884));
  XOR2_X1   g459(.A(G160), .B(new_n639), .Z(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(G162), .Z(new_n886));
  NAND3_X1  g461(.A1(new_n882), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(G37), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n886), .B1(new_n882), .B2(new_n884), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(KEYINPUT40), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n887), .A2(new_n888), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT40), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n893), .A2(new_n894), .A3(new_n890), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n892), .A2(new_n895), .ZN(G395));
  OR2_X1    g471(.A1(new_n611), .A2(G299), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n611), .A2(G299), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT41), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(KEYINPUT41), .A3(new_n898), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n625), .B(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n845), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n625), .B(KEYINPUT107), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n845), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n903), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n907), .A2(new_n909), .A3(new_n899), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT42), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n704), .B1(new_n589), .B2(new_n598), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n588), .A2(G305), .A3(new_n597), .A4(new_n595), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g490(.A(G303), .B(G288), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n913), .A2(new_n916), .A3(new_n914), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT42), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n907), .A2(new_n909), .A3(new_n899), .ZN(new_n923));
  AND2_X1   g498(.A1(new_n907), .A2(new_n909), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n922), .B(new_n923), .C1(new_n924), .C2(new_n903), .ZN(new_n925));
  AND3_X1   g500(.A1(new_n912), .A2(new_n921), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n921), .B1(new_n912), .B2(new_n925), .ZN(new_n927));
  OAI21_X1  g502(.A(G868), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(G868), .B2(new_n843), .ZN(G295));
  OAI21_X1  g504(.A(new_n928), .B1(G868), .B2(new_n843), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT110), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n913), .A2(new_n916), .A3(new_n914), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n916), .B1(new_n913), .B2(new_n914), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT109), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n918), .A2(new_n936), .A3(new_n919), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n566), .A2(G168), .A3(new_n568), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT108), .ZN(new_n940));
  NAND3_X1  g515(.A1(G171), .A2(new_n940), .A3(G286), .ZN(new_n941));
  OAI21_X1  g516(.A(KEYINPUT108), .B1(new_n540), .B2(G168), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n943), .A2(new_n845), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n845), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n898), .B(new_n897), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n906), .A2(new_n939), .A3(new_n941), .A4(new_n942), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n943), .A2(new_n845), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n901), .A2(new_n947), .A3(new_n902), .A4(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n938), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n932), .B1(new_n950), .B2(G37), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n899), .B1(new_n947), .B2(new_n948), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n944), .A2(new_n945), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n952), .B1(new_n903), .B2(new_n953), .ZN(new_n954));
  OAI211_X1 g529(.A(KEYINPUT110), .B(new_n888), .C1(new_n954), .C2(new_n938), .ZN(new_n955));
  AOI21_X1  g530(.A(KEYINPUT43), .B1(new_n954), .B2(new_n920), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n951), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n946), .A2(new_n949), .A3(new_n920), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n958), .B(new_n888), .C1(new_n954), .C2(new_n938), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT43), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n931), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT43), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  NOR3_X1   g538(.A1(new_n963), .A2(G37), .A3(new_n950), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n951), .A2(new_n955), .A3(new_n958), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n964), .B1(new_n965), .B2(KEYINPUT43), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n961), .B1(new_n931), .B2(new_n966), .ZN(G397));
  XOR2_X1   g542(.A(KEYINPUT111), .B(G1384), .Z(new_n968));
  NAND2_X1  g543(.A1(new_n878), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n471), .A2(new_n472), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(G2105), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(G40), .A3(new_n476), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n975), .A2(KEYINPUT112), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(KEYINPUT112), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n755), .B(G1996), .Z(new_n979));
  INV_X1    g554(.A(G2067), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n767), .B(new_n980), .ZN(new_n981));
  AND2_X1   g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  XNOR2_X1  g557(.A(new_n726), .B(new_n728), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n978), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n599), .A2(new_n717), .ZN(new_n985));
  NAND2_X1  g560(.A1(G290), .A2(G1986), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n978), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n984), .A2(new_n987), .ZN(new_n988));
  XOR2_X1   g563(.A(new_n988), .B(KEYINPUT113), .Z(new_n989));
  NAND2_X1  g564(.A1(G303), .A2(G8), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT55), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n990), .B(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT114), .ZN(new_n994));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n878), .A2(new_n994), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n491), .B1(new_n499), .B2(new_n496), .ZN(new_n997));
  OAI21_X1  g572(.A(KEYINPUT114), .B1(new_n997), .B2(G1384), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(new_n998), .A3(KEYINPUT50), .ZN(new_n999));
  INV_X1    g574(.A(G2090), .ZN(new_n1000));
  INV_X1    g575(.A(G40), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n473), .A2(new_n477), .A3(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n486), .A2(new_n493), .A3(new_n490), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n493), .B1(new_n486), .B2(new_n490), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n876), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1005), .A2(new_n1006), .A3(new_n995), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n999), .A2(new_n1000), .A3(new_n1002), .A4(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n878), .A2(KEYINPUT45), .A3(new_n968), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n1002), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT45), .B1(new_n1005), .B2(new_n995), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n701), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G8), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n993), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G1966), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n996), .A2(new_n998), .A3(new_n970), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1005), .A2(new_n995), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1002), .B1(new_n1018), .B2(new_n970), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1016), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n994), .B1(new_n878), .B2(new_n995), .ZN(new_n1021));
  NOR3_X1   g596(.A1(new_n997), .A2(KEYINPUT114), .A3(G1384), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1006), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n974), .B1(KEYINPUT50), .B2(new_n1018), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n1024), .A3(new_n793), .ZN(new_n1025));
  AOI211_X1 g600(.A(new_n1014), .B(G286), .C1(new_n1020), .C2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT49), .ZN(new_n1027));
  INV_X1    g602(.A(G1981), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n582), .A2(new_n583), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1028), .B1(new_n582), .B2(new_n583), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1027), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1002), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G305), .A2(G1981), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1034), .A2(KEYINPUT49), .A3(new_n1029), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1032), .A2(new_n1033), .A3(G8), .A4(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G288), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(G1976), .ZN(new_n1038));
  INV_X1    g613(.A(G1976), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT52), .B1(G288), .B2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1033), .A2(G8), .A3(new_n1038), .A4(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1036), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n996), .A2(new_n998), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1014), .B1(new_n1044), .B2(new_n1002), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1043), .B1(new_n1045), .B2(new_n1038), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1042), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(G164), .A2(G1384), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1002), .B1(new_n1048), .B2(new_n1006), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT50), .B1(new_n996), .B2(new_n998), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1049), .A2(new_n1050), .A3(G2090), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1012), .ZN(new_n1052));
  OAI211_X1 g627(.A(G8), .B(new_n992), .C1(new_n1051), .C2(new_n1052), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1015), .A2(new_n1026), .A3(new_n1047), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT63), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT117), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OR3_X1    g633(.A1(new_n1042), .A2(new_n1046), .A3(KEYINPUT115), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT115), .B1(new_n1042), .B2(new_n1046), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1053), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1062), .A2(new_n1055), .ZN(new_n1063));
  OAI21_X1  g638(.A(G8), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n993), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1061), .A2(new_n1063), .A3(new_n1026), .A4(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1054), .A2(KEYINPUT117), .A3(new_n1055), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1058), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n974), .B1(new_n996), .B2(new_n998), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1036), .A2(new_n1039), .A3(new_n1037), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1070), .A2(new_n1029), .ZN(new_n1071));
  AOI211_X1 g646(.A(new_n1014), .B(new_n1069), .C1(new_n1071), .C2(KEYINPUT116), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n1071), .A2(KEYINPUT116), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1072), .A2(new_n1073), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1015), .A2(new_n1047), .A3(new_n1053), .ZN(new_n1075));
  AND2_X1   g650(.A1(new_n1009), .A2(new_n1002), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1018), .A2(new_n970), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(new_n791), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G1961), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1076), .A2(KEYINPUT53), .A3(new_n791), .A4(new_n971), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1080), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT124), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT124), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1080), .A2(new_n1082), .A3(new_n1086), .A4(new_n1083), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(G171), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n974), .B1(new_n1048), .B2(KEYINPUT45), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n996), .A2(new_n998), .A3(new_n970), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1090), .A2(KEYINPUT53), .A3(new_n791), .A4(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1080), .A2(new_n1082), .A3(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1089), .B1(new_n1094), .B2(G301), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1075), .B1(new_n1088), .B2(new_n1095), .ZN(new_n1096));
  NOR3_X1   g671(.A1(new_n1049), .A2(new_n1050), .A3(G2084), .ZN(new_n1097));
  AOI21_X1  g672(.A(G1966), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1098));
  OAI21_X1  g673(.A(G8), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(G168), .A2(new_n1014), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(KEYINPUT51), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1099), .A2(KEYINPUT122), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1014), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1103));
  XOR2_X1   g678(.A(new_n1100), .B(KEYINPUT121), .Z(new_n1104));
  OAI21_X1  g679(.A(KEYINPUT51), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT122), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1101), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1106), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1102), .A2(new_n1105), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1100), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1093), .A2(new_n569), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1080), .A2(new_n1082), .A3(G301), .A4(new_n1083), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1112), .B1(new_n1115), .B2(new_n1089), .ZN(new_n1116));
  AOI211_X1 g691(.A(KEYINPUT123), .B(KEYINPUT54), .C1(new_n1113), .C2(new_n1114), .ZN(new_n1117));
  OAI211_X1 g692(.A(new_n1096), .B(new_n1111), .C1(new_n1116), .C2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1348), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1033), .B2(G2067), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1069), .A2(KEYINPUT118), .A3(new_n980), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1120), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n621), .ZN(new_n1125));
  XNOR2_X1  g700(.A(G299), .B(KEYINPUT57), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1007), .A2(new_n1002), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(G1956), .B1(new_n1128), .B2(new_n999), .ZN(new_n1129));
  XNOR2_X1  g704(.A(KEYINPUT56), .B(G2072), .ZN(new_n1130));
  AND4_X1   g705(.A1(new_n1002), .A2(new_n1077), .A3(new_n1009), .A4(new_n1130), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1126), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1125), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(G1956), .ZN(new_n1134));
  INV_X1    g709(.A(new_n999), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1134), .B1(new_n1135), .B2(new_n1127), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT57), .ZN(new_n1137));
  XNOR2_X1  g712(.A(G299), .B(new_n1137), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1076), .A2(new_n1077), .A3(new_n1130), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1136), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1133), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n1142));
  XOR2_X1   g717(.A(KEYINPUT119), .B(G1996), .Z(new_n1143));
  NAND3_X1  g718(.A1(new_n1076), .A2(new_n1077), .A3(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(KEYINPUT120), .B(KEYINPUT58), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(new_n810), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1033), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1142), .B1(new_n1148), .B2(new_n548), .ZN(new_n1149));
  AOI211_X1 g724(.A(KEYINPUT59), .B(new_n547), .C1(new_n1144), .C2(new_n1147), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1120), .A2(new_n1122), .A3(KEYINPUT60), .A4(new_n1123), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1149), .A2(new_n1150), .B1(new_n1151), .B2(new_n621), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1132), .A2(new_n1140), .A3(KEYINPUT61), .ZN(new_n1153));
  AOI21_X1  g728(.A(KEYINPUT61), .B1(new_n1132), .B2(new_n1140), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT60), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1124), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1157), .A2(new_n621), .A3(new_n1151), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1141), .B1(new_n1155), .B2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g734(.A(new_n1068), .B(new_n1074), .C1(new_n1118), .C2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1161), .B1(new_n1111), .B2(KEYINPUT62), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT62), .ZN(new_n1163));
  AOI211_X1 g738(.A(KEYINPUT125), .B(new_n1163), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1109), .A2(new_n1163), .A3(new_n1110), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1075), .A2(new_n1113), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g742(.A1(new_n1162), .A2(new_n1164), .A3(new_n1167), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n989), .B1(new_n1160), .B2(new_n1168), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT46), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1170), .B1(new_n978), .B2(G1996), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT126), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n869), .B(new_n981), .C1(new_n1170), .C2(G1996), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n976), .A2(new_n977), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1172), .A2(KEYINPUT47), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT48), .ZN(new_n1176));
  OR2_X1    g751(.A1(new_n978), .A2(new_n985), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n984), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1178), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1179));
  AND2_X1   g754(.A1(new_n867), .A2(new_n728), .ZN(new_n1180));
  AOI22_X1  g755(.A1(new_n982), .A2(new_n1180), .B1(new_n980), .B2(new_n768), .ZN(new_n1181));
  OAI211_X1 g756(.A(new_n1175), .B(new_n1179), .C1(new_n978), .C2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(KEYINPUT47), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1169), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  AND3_X1   g760(.A1(new_n672), .A2(G319), .A3(new_n657), .ZN(new_n1187));
  OAI21_X1  g761(.A(new_n1187), .B1(new_n695), .B2(new_n696), .ZN(new_n1188));
  NAND2_X1  g762(.A1(new_n1188), .A2(KEYINPUT127), .ZN(new_n1189));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n1190));
  OAI211_X1 g764(.A(new_n1187), .B(new_n1190), .C1(new_n695), .C2(new_n696), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n1189), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g766(.A(new_n1192), .B1(new_n893), .B2(new_n890), .ZN(new_n1193));
  NOR2_X1   g767(.A1(new_n1193), .A2(new_n966), .ZN(G308));
  NAND2_X1  g768(.A1(new_n965), .A2(KEYINPUT43), .ZN(new_n1195));
  INV_X1    g769(.A(new_n964), .ZN(new_n1196));
  NAND2_X1  g770(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n889), .A2(new_n891), .ZN(new_n1198));
  NAND3_X1  g772(.A1(new_n1197), .A2(new_n1198), .A3(new_n1192), .ZN(G225));
endmodule


