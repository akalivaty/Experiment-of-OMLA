

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579;

  AND2_X1 U320 ( .A1(G232GAT), .A2(G233GAT), .ZN(n288) );
  XNOR2_X1 U321 ( .A(n406), .B(n288), .ZN(n328) );
  NAND2_X1 U322 ( .A1(n536), .A2(n513), .ZN(n419) );
  XNOR2_X1 U323 ( .A(n329), .B(n328), .ZN(n331) );
  XNOR2_X1 U324 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U325 ( .A(n401), .B(KEYINPUT48), .ZN(n536) );
  XNOR2_X1 U326 ( .A(n339), .B(n338), .ZN(n344) );
  INV_X1 U327 ( .A(n536), .ZN(n539) );
  NOR2_X1 U328 ( .A1(n442), .A2(n522), .ZN(n556) );
  XOR2_X1 U329 ( .A(n441), .B(n440), .Z(n515) );
  XNOR2_X1 U330 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U331 ( .A(n446), .B(n445), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n423) );
  XNOR2_X1 U333 ( .A(G155GAT), .B(KEYINPUT87), .ZN(n289) );
  XNOR2_X1 U334 ( .A(n289), .B(KEYINPUT3), .ZN(n290) );
  XOR2_X1 U335 ( .A(n290), .B(KEYINPUT2), .Z(n292) );
  XNOR2_X1 U336 ( .A(G141GAT), .B(G162GAT), .ZN(n291) );
  XNOR2_X1 U337 ( .A(n292), .B(n291), .ZN(n317) );
  XOR2_X1 U338 ( .A(KEYINPUT86), .B(KEYINPUT21), .Z(n294) );
  XNOR2_X1 U339 ( .A(G218GAT), .B(KEYINPUT84), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U341 ( .A(n295), .B(KEYINPUT85), .Z(n297) );
  XNOR2_X1 U342 ( .A(G197GAT), .B(G211GAT), .ZN(n296) );
  XNOR2_X1 U343 ( .A(n297), .B(n296), .ZN(n418) );
  XNOR2_X1 U344 ( .A(n317), .B(n418), .ZN(n308) );
  XOR2_X1 U345 ( .A(KEYINPUT83), .B(G148GAT), .Z(n299) );
  XNOR2_X1 U346 ( .A(G50GAT), .B(G22GAT), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n301) );
  XNOR2_X1 U348 ( .A(G106GAT), .B(G78GAT), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n300), .B(G204GAT), .ZN(n387) );
  XOR2_X1 U350 ( .A(n301), .B(n387), .Z(n306) );
  XOR2_X1 U351 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n303) );
  NAND2_X1 U352 ( .A1(G228GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U353 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U354 ( .A(KEYINPUT22), .B(n304), .ZN(n305) );
  XNOR2_X1 U355 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n465) );
  XOR2_X1 U357 ( .A(G127GAT), .B(KEYINPUT79), .Z(n310) );
  XNOR2_X1 U358 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n430) );
  XNOR2_X1 U360 ( .A(G120GAT), .B(G148GAT), .ZN(n311) );
  XNOR2_X1 U361 ( .A(n311), .B(G57GAT), .ZN(n375) );
  XNOR2_X1 U362 ( .A(n430), .B(n375), .ZN(n325) );
  XOR2_X1 U363 ( .A(KEYINPUT1), .B(KEYINPUT88), .Z(n313) );
  XNOR2_X1 U364 ( .A(KEYINPUT5), .B(KEYINPUT4), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n315) );
  XOR2_X1 U366 ( .A(G1GAT), .B(G85GAT), .Z(n314) );
  XNOR2_X1 U367 ( .A(n315), .B(n314), .ZN(n321) );
  XOR2_X1 U368 ( .A(KEYINPUT6), .B(KEYINPUT89), .Z(n319) );
  XNOR2_X1 U369 ( .A(G29GAT), .B(G134GAT), .ZN(n316) );
  XNOR2_X1 U370 ( .A(n316), .B(KEYINPUT76), .ZN(n342) );
  XNOR2_X1 U371 ( .A(n317), .B(n342), .ZN(n318) );
  XNOR2_X1 U372 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n323) );
  NAND2_X1 U374 ( .A1(G225GAT), .A2(G233GAT), .ZN(n322) );
  XNOR2_X1 U375 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U376 ( .A(n325), .B(n324), .ZN(n463) );
  XNOR2_X1 U377 ( .A(KEYINPUT90), .B(n463), .ZN(n510) );
  INV_X1 U378 ( .A(n510), .ZN(n558) );
  AND2_X1 U379 ( .A1(n465), .A2(n558), .ZN(n421) );
  XOR2_X1 U380 ( .A(KEYINPUT54), .B(KEYINPUT119), .Z(n420) );
  XOR2_X1 U381 ( .A(KEYINPUT65), .B(G106GAT), .Z(n327) );
  XNOR2_X1 U382 ( .A(G162GAT), .B(G218GAT), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n327), .B(n326), .ZN(n329) );
  XOR2_X1 U384 ( .A(G36GAT), .B(G190GAT), .Z(n406) );
  INV_X1 U385 ( .A(KEYINPUT75), .ZN(n330) );
  XNOR2_X1 U386 ( .A(n331), .B(n330), .ZN(n339) );
  XOR2_X1 U387 ( .A(G43GAT), .B(G50GAT), .Z(n333) );
  XNOR2_X1 U388 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n372) );
  XNOR2_X1 U390 ( .A(n372), .B(KEYINPUT74), .ZN(n337) );
  XOR2_X1 U391 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n335) );
  XNOR2_X1 U392 ( .A(KEYINPUT73), .B(KEYINPUT10), .ZN(n334) );
  XOR2_X1 U393 ( .A(n335), .B(n334), .Z(n336) );
  XOR2_X1 U394 ( .A(G85GAT), .B(KEYINPUT70), .Z(n341) );
  XNOR2_X1 U395 ( .A(G99GAT), .B(G92GAT), .ZN(n340) );
  XNOR2_X1 U396 ( .A(n341), .B(n340), .ZN(n386) );
  XNOR2_X1 U397 ( .A(n386), .B(n342), .ZN(n343) );
  XOR2_X1 U398 ( .A(n344), .B(n343), .Z(n550) );
  INV_X1 U399 ( .A(n550), .ZN(n450) );
  XOR2_X1 U400 ( .A(G8GAT), .B(G183GAT), .Z(n402) );
  XNOR2_X1 U401 ( .A(G22GAT), .B(G15GAT), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n345), .B(G1GAT), .ZN(n359) );
  XOR2_X1 U403 ( .A(n402), .B(n359), .Z(n347) );
  NAND2_X1 U404 ( .A1(G231GAT), .A2(G233GAT), .ZN(n346) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U406 ( .A(G71GAT), .B(KEYINPUT13), .Z(n378) );
  XOR2_X1 U407 ( .A(n348), .B(n378), .Z(n350) );
  XNOR2_X1 U408 ( .A(G155GAT), .B(G78GAT), .ZN(n349) );
  XNOR2_X1 U409 ( .A(n350), .B(n349), .ZN(n358) );
  XOR2_X1 U410 ( .A(G57GAT), .B(G64GAT), .Z(n352) );
  XNOR2_X1 U411 ( .A(G127GAT), .B(G211GAT), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U413 ( .A(KEYINPUT15), .B(KEYINPUT77), .Z(n354) );
  XNOR2_X1 U414 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n353) );
  XNOR2_X1 U415 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U416 ( .A(n356), .B(n355), .Z(n357) );
  XOR2_X1 U417 ( .A(n358), .B(n357), .Z(n555) );
  INV_X1 U418 ( .A(n555), .ZN(n571) );
  NAND2_X1 U419 ( .A1(n450), .A2(n571), .ZN(n393) );
  XOR2_X1 U420 ( .A(KEYINPUT110), .B(KEYINPUT46), .Z(n391) );
  XOR2_X1 U421 ( .A(G29GAT), .B(n359), .Z(n361) );
  NAND2_X1 U422 ( .A1(G229GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U423 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U424 ( .A(n362), .B(G36GAT), .Z(n370) );
  XOR2_X1 U425 ( .A(G113GAT), .B(G197GAT), .Z(n364) );
  XNOR2_X1 U426 ( .A(G169GAT), .B(G141GAT), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U428 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n366) );
  XNOR2_X1 U429 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U431 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U433 ( .A(n371), .B(KEYINPUT66), .Z(n374) );
  XNOR2_X1 U434 ( .A(n372), .B(KEYINPUT67), .ZN(n373) );
  XOR2_X1 U435 ( .A(n374), .B(n373), .Z(n562) );
  INV_X1 U436 ( .A(n562), .ZN(n552) );
  XOR2_X1 U437 ( .A(G176GAT), .B(G64GAT), .Z(n403) );
  XOR2_X1 U438 ( .A(n375), .B(n403), .Z(n377) );
  NAND2_X1 U439 ( .A1(G230GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U440 ( .A(n377), .B(n376), .ZN(n379) );
  XOR2_X1 U441 ( .A(n379), .B(n378), .Z(n381) );
  XNOR2_X1 U442 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U444 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n383) );
  XNOR2_X1 U445 ( .A(KEYINPUT31), .B(KEYINPUT69), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U447 ( .A(n385), .B(n384), .Z(n389) );
  XNOR2_X1 U448 ( .A(n387), .B(n386), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n567) );
  XNOR2_X1 U450 ( .A(n567), .B(KEYINPUT41), .ZN(n541) );
  NAND2_X1 U451 ( .A1(n552), .A2(n541), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n391), .B(n390), .ZN(n392) );
  NOR2_X1 U453 ( .A1(n393), .A2(n392), .ZN(n394) );
  XNOR2_X1 U454 ( .A(KEYINPUT47), .B(n394), .ZN(n400) );
  XOR2_X1 U455 ( .A(KEYINPUT36), .B(n550), .Z(n577) );
  NOR2_X1 U456 ( .A1(n577), .A2(n571), .ZN(n395) );
  XNOR2_X1 U457 ( .A(KEYINPUT45), .B(n395), .ZN(n396) );
  NAND2_X1 U458 ( .A1(n396), .A2(n567), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n397), .B(KEYINPUT111), .ZN(n398) );
  NAND2_X1 U460 ( .A1(n398), .A2(n562), .ZN(n399) );
  NAND2_X1 U461 ( .A1(n400), .A2(n399), .ZN(n401) );
  XOR2_X1 U462 ( .A(n403), .B(n402), .Z(n405) );
  NAND2_X1 U463 ( .A1(G226GAT), .A2(G233GAT), .ZN(n404) );
  XNOR2_X1 U464 ( .A(n405), .B(n404), .ZN(n407) );
  XOR2_X1 U465 ( .A(n407), .B(n406), .Z(n416) );
  XOR2_X1 U466 ( .A(KEYINPUT94), .B(KEYINPUT91), .Z(n409) );
  XNOR2_X1 U467 ( .A(G204GAT), .B(G92GAT), .ZN(n408) );
  XNOR2_X1 U468 ( .A(n409), .B(n408), .ZN(n414) );
  XOR2_X1 U469 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n411) );
  XNOR2_X1 U470 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n410) );
  XNOR2_X1 U471 ( .A(n411), .B(n410), .ZN(n431) );
  XNOR2_X1 U472 ( .A(n431), .B(KEYINPUT92), .ZN(n412) );
  XNOR2_X1 U473 ( .A(n412), .B(KEYINPUT93), .ZN(n413) );
  XNOR2_X1 U474 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U475 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n513) );
  XOR2_X1 U477 ( .A(n420), .B(n419), .Z(n559) );
  NAND2_X1 U478 ( .A1(n421), .A2(n559), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n442) );
  XOR2_X1 U480 ( .A(KEYINPUT20), .B(G183GAT), .Z(n425) );
  XNOR2_X1 U481 ( .A(G176GAT), .B(G120GAT), .ZN(n424) );
  XNOR2_X1 U482 ( .A(n425), .B(n424), .ZN(n441) );
  XOR2_X1 U483 ( .A(KEYINPUT64), .B(G71GAT), .Z(n427) );
  XNOR2_X1 U484 ( .A(G190GAT), .B(G134GAT), .ZN(n426) );
  XNOR2_X1 U485 ( .A(n427), .B(n426), .ZN(n429) );
  XOR2_X1 U486 ( .A(G43GAT), .B(G99GAT), .Z(n428) );
  XNOR2_X1 U487 ( .A(n429), .B(n428), .ZN(n437) );
  XNOR2_X1 U488 ( .A(n431), .B(n430), .ZN(n435) );
  XOR2_X1 U489 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n433) );
  XNOR2_X1 U490 ( .A(G15GAT), .B(KEYINPUT80), .ZN(n432) );
  XNOR2_X1 U491 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n439) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U495 ( .A(n439), .B(n438), .ZN(n440) );
  INV_X1 U496 ( .A(n515), .ZN(n522) );
  NAND2_X1 U497 ( .A1(n556), .A2(n550), .ZN(n446) );
  XOR2_X1 U498 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n444) );
  INV_X1 U499 ( .A(G190GAT), .ZN(n443) );
  NAND2_X1 U500 ( .A1(n556), .A2(n541), .ZN(n449) );
  XOR2_X1 U501 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n447) );
  XNOR2_X1 U502 ( .A(n447), .B(G176GAT), .ZN(n448) );
  XNOR2_X1 U503 ( .A(n449), .B(n448), .ZN(G1349GAT) );
  XNOR2_X1 U504 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n473) );
  NAND2_X1 U505 ( .A1(n552), .A2(n567), .ZN(n484) );
  XOR2_X1 U506 ( .A(KEYINPUT78), .B(KEYINPUT16), .Z(n452) );
  NAND2_X1 U507 ( .A1(n555), .A2(n450), .ZN(n451) );
  XNOR2_X1 U508 ( .A(n452), .B(n451), .ZN(n470) );
  NAND2_X1 U509 ( .A1(n515), .A2(n513), .ZN(n453) );
  XNOR2_X1 U510 ( .A(KEYINPUT98), .B(n453), .ZN(n454) );
  NAND2_X1 U511 ( .A1(n454), .A2(n465), .ZN(n455) );
  XNOR2_X1 U512 ( .A(KEYINPUT25), .B(n455), .ZN(n461) );
  XNOR2_X1 U513 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n457) );
  NOR2_X1 U514 ( .A1(n515), .A2(n465), .ZN(n456) );
  XNOR2_X1 U515 ( .A(n457), .B(n456), .ZN(n560) );
  XOR2_X1 U516 ( .A(KEYINPUT27), .B(KEYINPUT95), .Z(n458) );
  XNOR2_X1 U517 ( .A(n513), .B(n458), .ZN(n464) );
  NAND2_X1 U518 ( .A1(n560), .A2(n464), .ZN(n459) );
  XNOR2_X1 U519 ( .A(KEYINPUT97), .B(n459), .ZN(n460) );
  NOR2_X1 U520 ( .A1(n461), .A2(n460), .ZN(n462) );
  NOR2_X1 U521 ( .A1(n463), .A2(n462), .ZN(n468) );
  AND2_X1 U522 ( .A1(n510), .A2(n464), .ZN(n537) );
  XOR2_X1 U523 ( .A(n465), .B(KEYINPUT28), .Z(n517) );
  INV_X1 U524 ( .A(n517), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n537), .A2(n466), .ZN(n521) );
  NOR2_X1 U526 ( .A1(n515), .A2(n521), .ZN(n467) );
  NOR2_X1 U527 ( .A1(n468), .A2(n467), .ZN(n481) );
  INV_X1 U528 ( .A(n481), .ZN(n469) );
  NAND2_X1 U529 ( .A1(n470), .A2(n469), .ZN(n499) );
  NOR2_X1 U530 ( .A1(n484), .A2(n499), .ZN(n471) );
  XOR2_X1 U531 ( .A(KEYINPUT99), .B(n471), .Z(n479) );
  NAND2_X1 U532 ( .A1(n479), .A2(n510), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n473), .B(n472), .ZN(G1324GAT) );
  NAND2_X1 U534 ( .A1(n513), .A2(n479), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n474), .B(KEYINPUT100), .ZN(n475) );
  XNOR2_X1 U536 ( .A(G8GAT), .B(n475), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n477) );
  NAND2_X1 U538 ( .A1(n479), .A2(n515), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U540 ( .A(G15GAT), .B(n478), .Z(G1326GAT) );
  NAND2_X1 U541 ( .A1(n479), .A2(n517), .ZN(n480) );
  XNOR2_X1 U542 ( .A(n480), .B(G22GAT), .ZN(G1327GAT) );
  NOR2_X1 U543 ( .A1(n481), .A2(n577), .ZN(n482) );
  NAND2_X1 U544 ( .A1(n571), .A2(n482), .ZN(n483) );
  XOR2_X1 U545 ( .A(KEYINPUT37), .B(n483), .Z(n509) );
  NOR2_X1 U546 ( .A1(n509), .A2(n484), .ZN(n486) );
  XNOR2_X1 U547 ( .A(KEYINPUT38), .B(KEYINPUT102), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n495) );
  NAND2_X1 U549 ( .A1(n495), .A2(n510), .ZN(n488) );
  XOR2_X1 U550 ( .A(G29GAT), .B(KEYINPUT39), .Z(n487) );
  XNOR2_X1 U551 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  XOR2_X1 U552 ( .A(G36GAT), .B(KEYINPUT103), .Z(n490) );
  NAND2_X1 U553 ( .A1(n495), .A2(n513), .ZN(n489) );
  XNOR2_X1 U554 ( .A(n490), .B(n489), .ZN(G1329GAT) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(KEYINPUT104), .ZN(n494) );
  XOR2_X1 U556 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n492) );
  NAND2_X1 U557 ( .A1(n495), .A2(n515), .ZN(n491) );
  XNOR2_X1 U558 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U559 ( .A(n494), .B(n493), .ZN(G1330GAT) );
  NAND2_X1 U560 ( .A1(n495), .A2(n517), .ZN(n496) );
  XNOR2_X1 U561 ( .A(n496), .B(KEYINPUT106), .ZN(n497) );
  XNOR2_X1 U562 ( .A(G50GAT), .B(n497), .ZN(G1331GAT) );
  XOR2_X1 U563 ( .A(KEYINPUT42), .B(KEYINPUT108), .Z(n501) );
  NAND2_X1 U564 ( .A1(n541), .A2(n562), .ZN(n498) );
  XOR2_X1 U565 ( .A(KEYINPUT107), .B(n498), .Z(n508) );
  NOR2_X1 U566 ( .A1(n499), .A2(n508), .ZN(n505) );
  NAND2_X1 U567 ( .A1(n505), .A2(n510), .ZN(n500) );
  XNOR2_X1 U568 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U569 ( .A(G57GAT), .B(n502), .Z(G1332GAT) );
  NAND2_X1 U570 ( .A1(n513), .A2(n505), .ZN(n503) );
  XNOR2_X1 U571 ( .A(n503), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n505), .A2(n515), .ZN(n504) );
  XNOR2_X1 U573 ( .A(n504), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .Z(n507) );
  NAND2_X1 U575 ( .A1(n505), .A2(n517), .ZN(n506) );
  XNOR2_X1 U576 ( .A(n507), .B(n506), .ZN(G1335GAT) );
  XOR2_X1 U577 ( .A(G85GAT), .B(KEYINPUT109), .Z(n512) );
  NOR2_X1 U578 ( .A1(n509), .A2(n508), .ZN(n518) );
  NAND2_X1 U579 ( .A1(n518), .A2(n510), .ZN(n511) );
  XNOR2_X1 U580 ( .A(n512), .B(n511), .ZN(G1336GAT) );
  NAND2_X1 U581 ( .A1(n513), .A2(n518), .ZN(n514) );
  XNOR2_X1 U582 ( .A(n514), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U583 ( .A1(n518), .A2(n515), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n516), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U585 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n519), .B(KEYINPUT44), .ZN(n520) );
  XNOR2_X1 U587 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  NOR2_X1 U588 ( .A1(n522), .A2(n521), .ZN(n523) );
  NAND2_X1 U589 ( .A1(n523), .A2(n536), .ZN(n524) );
  XOR2_X1 U590 ( .A(KEYINPUT112), .B(n524), .Z(n532) );
  NAND2_X1 U591 ( .A1(n532), .A2(n552), .ZN(n525) );
  XNOR2_X1 U592 ( .A(n525), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(G120GAT), .B(KEYINPUT49), .Z(n527) );
  NAND2_X1 U594 ( .A1(n532), .A2(n541), .ZN(n526) );
  XNOR2_X1 U595 ( .A(n527), .B(n526), .ZN(G1341GAT) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n531) );
  XOR2_X1 U597 ( .A(KEYINPUT114), .B(KEYINPUT113), .Z(n529) );
  NAND2_X1 U598 ( .A1(n555), .A2(n532), .ZN(n528) );
  XNOR2_X1 U599 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U600 ( .A(n531), .B(n530), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n534) );
  NAND2_X1 U602 ( .A1(n532), .A2(n550), .ZN(n533) );
  XNOR2_X1 U603 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U604 ( .A(G134GAT), .B(n535), .Z(G1343GAT) );
  NAND2_X1 U605 ( .A1(n560), .A2(n537), .ZN(n538) );
  NOR2_X1 U606 ( .A1(n539), .A2(n538), .ZN(n549) );
  NAND2_X1 U607 ( .A1(n552), .A2(n549), .ZN(n540) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(n540), .ZN(G1344GAT) );
  NAND2_X1 U609 ( .A1(n541), .A2(n549), .ZN(n547) );
  XOR2_X1 U610 ( .A(KEYINPUT118), .B(KEYINPUT117), .Z(n543) );
  XNOR2_X1 U611 ( .A(KEYINPUT116), .B(KEYINPUT53), .ZN(n542) );
  XNOR2_X1 U612 ( .A(n543), .B(n542), .ZN(n545) );
  XOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT52), .Z(n544) );
  XNOR2_X1 U614 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(G1345GAT) );
  NAND2_X1 U616 ( .A1(n549), .A2(n555), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n548), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n551), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n552), .A2(n556), .ZN(n554) );
  XOR2_X1 U621 ( .A(G169GAT), .B(KEYINPUT121), .Z(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(G1348GAT) );
  NAND2_X1 U623 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(G183GAT), .ZN(G1350GAT) );
  AND2_X1 U625 ( .A1(n559), .A2(n558), .ZN(n561) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n576) );
  NOR2_X1 U627 ( .A1(n576), .A2(n562), .ZN(n566) );
  XOR2_X1 U628 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n564) );
  XNOR2_X1 U629 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(G1352GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n576), .ZN(n569) );
  XNOR2_X1 U633 ( .A(KEYINPUT124), .B(KEYINPUT61), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G204GAT), .B(n570), .ZN(G1353GAT) );
  NOR2_X1 U636 ( .A1(n571), .A2(n576), .ZN(n573) );
  XNOR2_X1 U637 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n573), .B(n572), .ZN(G1354GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n575) );
  XNOR2_X1 U640 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n579) );
  NOR2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(n579), .B(n578), .Z(G1355GAT) );
endmodule

