//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:33 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n730, new_n731, new_n732, new_n733, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003;
  INV_X1    g000(.A(KEYINPUT98), .ZN(new_n202));
  INV_X1    g001(.A(G57gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G64gat), .ZN(new_n204));
  INV_X1    g003(.A(G64gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G57gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT9), .ZN(new_n207));
  NAND2_X1  g006(.A1(G71gat), .A2(G78gat), .ZN(new_n208));
  AOI22_X1  g007(.A1(new_n204), .A2(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  OR2_X1    g008(.A1(G71gat), .A2(G78gat), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n210), .A2(KEYINPUT97), .A3(new_n208), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT97), .B1(new_n210), .B2(new_n208), .ZN(new_n213));
  OAI211_X1 g012(.A(new_n202), .B(new_n209), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n204), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n208), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n213), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n217), .B1(new_n218), .B2(new_n211), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n210), .A2(new_n208), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT98), .B1(new_n209), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n214), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT21), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G231gat), .A2(G233gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(G127gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(G183gat), .B(G211gat), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XOR2_X1   g029(.A(G15gat), .B(G22gat), .Z(new_n231));
  INV_X1    g030(.A(G1gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G15gat), .B(G22gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT16), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n234), .B1(new_n235), .B2(G1gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n233), .A2(new_n236), .A3(KEYINPUT92), .ZN(new_n237));
  INV_X1    g036(.A(G8gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT94), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n237), .B(G8gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT94), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n240), .B(new_n243), .C1(new_n224), .C2(new_n223), .ZN(new_n244));
  XNOR2_X1  g043(.A(new_n244), .B(KEYINPUT99), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n246));
  INV_X1    g045(.A(G155gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n245), .B(new_n248), .Z(new_n249));
  OR2_X1    g048(.A1(new_n230), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n249), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  OR2_X1    g051(.A1(KEYINPUT101), .A2(G92gat), .ZN(new_n253));
  INV_X1    g052(.A(G85gat), .ZN(new_n254));
  NAND2_X1  g053(.A1(KEYINPUT101), .A2(G92gat), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G99gat), .ZN(new_n257));
  INV_X1    g056(.A(G106gat), .ZN(new_n258));
  OAI21_X1  g057(.A(KEYINPUT8), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G99gat), .B(G106gat), .Z(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G85gat), .A2(G92gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(KEYINPUT100), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT100), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n265), .A2(G85gat), .A3(G92gat), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT7), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n264), .A2(new_n266), .A3(KEYINPUT7), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n260), .A2(new_n262), .A3(new_n268), .A4(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n269), .A2(new_n259), .A3(new_n256), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n261), .B1(new_n271), .B2(new_n267), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n270), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G36gat), .ZN(new_n274));
  AND2_X1   g073(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G29gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n278), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n280), .A2(KEYINPUT15), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(KEYINPUT15), .ZN(new_n282));
  XNOR2_X1  g081(.A(G43gat), .B(G50gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n282), .A2(new_n283), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(KEYINPUT17), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT17), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n288), .B1(new_n284), .B2(new_n285), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n273), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  AND3_X1   g089(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n273), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n291), .B1(new_n286), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  XNOR2_X1  g093(.A(G190gat), .B(G218gat), .ZN(new_n295));
  XNOR2_X1  g094(.A(new_n295), .B(KEYINPUT102), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n294), .B(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT103), .ZN(new_n299));
  INV_X1    g098(.A(new_n296), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n299), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT104), .ZN(new_n302));
  XNOR2_X1  g101(.A(G134gat), .B(G162gat), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n301), .A2(new_n302), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n302), .B1(new_n301), .B2(new_n305), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n298), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n308), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n310), .A2(new_n297), .A3(new_n306), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n252), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT106), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT10), .ZN(new_n316));
  NOR3_X1   g115(.A1(new_n223), .A2(new_n273), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n270), .A2(KEYINPUT105), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n222), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(new_n292), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n273), .A2(new_n318), .A3(new_n222), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n317), .B1(new_n322), .B2(new_n316), .ZN(new_n323));
  NAND2_X1  g122(.A1(G230gat), .A2(G233gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n315), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT10), .B1(new_n320), .B2(new_n321), .ZN(new_n327));
  OAI211_X1 g126(.A(KEYINPUT106), .B(new_n324), .C1(new_n327), .C2(new_n317), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n320), .A2(new_n325), .A3(new_n321), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  XNOR2_X1  g130(.A(G120gat), .B(G148gat), .ZN(new_n332));
  XNOR2_X1  g131(.A(G176gat), .B(G204gat), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n332), .B(new_n333), .Z(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n329), .A2(new_n336), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n323), .A2(new_n325), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n335), .B1(new_n338), .B2(new_n331), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n314), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G78gat), .B(G106gat), .ZN(new_n342));
  XNOR2_X1  g141(.A(KEYINPUT31), .B(G50gat), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n342), .B(new_n343), .Z(new_n344));
  NAND2_X1  g143(.A1(G228gat), .A2(G233gat), .ZN(new_n345));
  INV_X1    g144(.A(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G148gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT75), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G148gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n350), .A3(G141gat), .ZN(new_n351));
  OR2_X1    g150(.A1(new_n347), .A2(G141gat), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT76), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n351), .A2(KEYINPUT76), .A3(new_n352), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n357));
  AND2_X1   g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(G155gat), .A2(G162gat), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G162gat), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n247), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G155gat), .A2(G162gat), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n362), .A2(KEYINPUT77), .A3(new_n363), .ZN(new_n364));
  AOI22_X1  g163(.A1(new_n360), .A2(new_n364), .B1(KEYINPUT2), .B2(new_n363), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n355), .A2(new_n356), .A3(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G141gat), .B(G148gat), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n363), .B(new_n362), .C1(new_n367), .C2(KEYINPUT2), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G197gat), .B(G204gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT73), .B(G211gat), .ZN(new_n371));
  INV_X1    g170(.A(G218gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n370), .B1(new_n373), .B2(KEYINPUT22), .ZN(new_n374));
  XNOR2_X1  g173(.A(G211gat), .B(G218gat), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n370), .B(new_n375), .C1(new_n373), .C2(KEYINPUT22), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT29), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n369), .B1(new_n379), .B2(KEYINPUT3), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT84), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(new_n378), .ZN(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT3), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n366), .A2(new_n384), .A3(new_n368), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n380), .A2(new_n381), .B1(new_n383), .B2(new_n387), .ZN(new_n388));
  OAI211_X1 g187(.A(KEYINPUT84), .B(new_n369), .C1(new_n379), .C2(KEYINPUT3), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n346), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n380), .A2(new_n346), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n385), .A2(new_n392), .A3(new_n386), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n382), .B1(new_n387), .B2(KEYINPUT85), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n391), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT86), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n344), .B1(new_n396), .B2(G22gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n380), .A2(new_n381), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n387), .A2(new_n383), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n389), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n345), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT86), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n394), .A2(new_n393), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n404), .A2(new_n346), .A3(new_n380), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n402), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n396), .A2(new_n406), .A3(G22gat), .ZN(new_n407));
  NAND2_X1  g206(.A1(KEYINPUT87), .A2(G22gat), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n402), .A2(new_n405), .A3(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n344), .ZN(new_n410));
  AND2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI211_X1 g210(.A(KEYINPUT87), .B(G22gat), .C1(new_n390), .C2(new_n395), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n398), .A2(new_n407), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(G1gat), .B(G29gat), .Z(new_n414));
  XNOR2_X1  g213(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G57gat), .B(G85gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G120gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(G113gat), .ZN(new_n421));
  INV_X1    g220(.A(G113gat), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G120gat), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT1), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G134gat), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n425), .A2(G127gat), .ZN(new_n426));
  INV_X1    g225(.A(G127gat), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n427), .A2(G134gat), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT69), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT69), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n430), .B1(new_n425), .B2(G127gat), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n424), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n426), .A2(new_n428), .ZN(new_n433));
  AND2_X1   g232(.A1(new_n433), .A2(new_n424), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n435), .A2(new_n366), .A3(new_n368), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT4), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT4), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n435), .A2(new_n366), .A3(new_n438), .A4(new_n368), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n369), .A2(KEYINPUT3), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n433), .A2(new_n424), .ZN(new_n442));
  INV_X1    g241(.A(new_n431), .ZN(new_n443));
  XOR2_X1   g242(.A(G127gat), .B(G134gat), .Z(new_n444));
  AOI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(KEYINPUT69), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n442), .B1(new_n445), .B2(new_n424), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n441), .A2(new_n446), .A3(new_n385), .ZN(new_n447));
  XOR2_X1   g246(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(G225gat), .A2(G233gat), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n440), .A2(new_n447), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT82), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n440), .A2(new_n447), .A3(KEYINPUT82), .A4(new_n452), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n437), .A2(KEYINPUT78), .A3(new_n439), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT78), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n436), .A2(new_n459), .A3(KEYINPUT4), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n458), .A2(new_n447), .A3(new_n450), .A4(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT80), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n369), .A2(new_n446), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n450), .B1(new_n463), .B2(new_n436), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n464), .B2(new_n448), .ZN(new_n465));
  INV_X1    g264(.A(new_n436), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n435), .B1(new_n368), .B2(new_n366), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n451), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n468), .A2(KEYINPUT80), .A3(new_n449), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n461), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n419), .B1(new_n457), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT6), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT6), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n457), .A2(new_n470), .A3(new_n419), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT83), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n473), .B(new_n474), .C1(new_n471), .C2(new_n475), .ZN(new_n476));
  AND2_X1   g275(.A1(new_n471), .A2(new_n475), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n472), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(G8gat), .B(G36gat), .ZN(new_n479));
  XNOR2_X1  g278(.A(G64gat), .B(G92gat), .ZN(new_n480));
  XOR2_X1   g279(.A(new_n479), .B(new_n480), .Z(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  AND2_X1   g281(.A1(G226gat), .A2(G233gat), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n483), .A2(KEYINPUT29), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n486));
  INV_X1    g285(.A(G169gat), .ZN(new_n487));
  INV_X1    g286(.A(G176gat), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT23), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT24), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n490), .A2(G183gat), .A3(G190gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(G169gat), .A2(G176gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(G183gat), .A2(G190gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT24), .ZN(new_n495));
  NOR2_X1   g294(.A1(G183gat), .A2(G190gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(G169gat), .A2(G176gat), .ZN(new_n499));
  OAI21_X1  g298(.A(KEYINPUT65), .B1(new_n499), .B2(KEYINPUT23), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT65), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT23), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n501), .B(new_n502), .C1(G169gat), .C2(G176gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n486), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT25), .ZN(new_n506));
  AND3_X1   g305(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n495), .A2(new_n496), .ZN(new_n508));
  AND4_X1   g307(.A1(new_n506), .A2(new_n507), .A3(new_n504), .A4(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT26), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT26), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(G169gat), .B2(G176gat), .ZN(new_n513));
  AND2_X1   g312(.A1(G169gat), .A2(G176gat), .ZN(new_n514));
  OAI211_X1 g313(.A(new_n511), .B(new_n494), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT68), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n487), .A2(new_n488), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n518), .A2(new_n512), .A3(new_n492), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n519), .A2(KEYINPUT68), .A3(new_n494), .A4(new_n511), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT27), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G183gat), .ZN(new_n522));
  INV_X1    g321(.A(G183gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT27), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT28), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n526), .A2(G190gat), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  OAI21_X1  g327(.A(KEYINPUT67), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT27), .B(G183gat), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT67), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(new_n531), .A3(new_n527), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n525), .A2(KEYINPUT66), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT66), .ZN(new_n535));
  AOI21_X1  g334(.A(G190gat), .B1(new_n522), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(KEYINPUT28), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  OAI211_X1 g336(.A(new_n517), .B(new_n520), .C1(new_n533), .C2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n485), .B1(new_n510), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n517), .A2(new_n520), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n529), .A2(new_n532), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n534), .A2(new_n536), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n526), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n540), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n507), .A2(new_n504), .A3(new_n508), .ZN(new_n545));
  INV_X1    g344(.A(new_n486), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n498), .A2(new_n506), .A3(new_n504), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g348(.A(KEYINPUT74), .B1(new_n544), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT74), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n510), .A2(new_n551), .A3(new_n538), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n539), .B1(new_n553), .B2(new_n483), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n554), .A2(new_n383), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n550), .A2(new_n552), .A3(new_n484), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n510), .A2(new_n483), .A3(new_n538), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n556), .A2(new_n383), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n482), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n558), .B(new_n481), .C1(new_n554), .C2(new_n383), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(KEYINPUT30), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n558), .B1(new_n554), .B2(new_n383), .ZN(new_n563));
  OR3_X1    g362(.A1(new_n563), .A2(KEYINPUT30), .A3(new_n482), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n478), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT34), .ZN(new_n567));
  OAI211_X1 g366(.A(KEYINPUT70), .B(new_n435), .C1(new_n544), .C2(new_n549), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n435), .A2(KEYINPUT70), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT70), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n446), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n510), .A2(new_n569), .A3(new_n538), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G227gat), .ZN(new_n574));
  INV_X1    g373(.A(G233gat), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n567), .B1(new_n573), .B2(new_n577), .ZN(new_n578));
  AOI211_X1 g377(.A(KEYINPUT34), .B(new_n576), .C1(new_n568), .C2(new_n572), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n568), .A2(new_n572), .A3(new_n576), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT32), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT33), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G15gat), .B(G43gat), .Z(new_n585));
  XNOR2_X1  g384(.A(G71gat), .B(G99gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n582), .A2(new_n584), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n587), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n581), .B(KEYINPUT32), .C1(new_n583), .C2(new_n589), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n580), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n578), .ZN(new_n592));
  INV_X1    g391(.A(new_n579), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n588), .A2(new_n590), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT72), .B1(new_n591), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n588), .A2(new_n590), .ZN(new_n596));
  INV_X1    g395(.A(new_n580), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n588), .A3(new_n590), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(KEYINPUT71), .A3(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT71), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n594), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n595), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(KEYINPUT36), .ZN(new_n604));
  AOI211_X1 g403(.A(KEYINPUT72), .B(KEYINPUT36), .C1(new_n598), .C2(new_n599), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n413), .A2(new_n566), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n474), .A2(new_n473), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n472), .B1(new_n608), .B2(new_n471), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT38), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n554), .A2(new_n382), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n556), .A2(new_n382), .A3(new_n557), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT37), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n610), .B1(new_n611), .B2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(KEYINPUT89), .B(KEYINPUT37), .Z(new_n615));
  OAI211_X1 g414(.A(new_n558), .B(new_n615), .C1(new_n554), .C2(new_n383), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n482), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n561), .B1(new_n614), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(KEYINPUT90), .B1(new_n609), .B2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n561), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n616), .A2(new_n482), .ZN(new_n621));
  AND2_X1   g420(.A1(new_n612), .A2(KEYINPUT37), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n553), .A2(new_n483), .ZN(new_n623));
  OAI21_X1  g422(.A(new_n383), .B1(new_n623), .B2(new_n539), .ZN(new_n624));
  AOI21_X1  g423(.A(KEYINPUT38), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n620), .B1(new_n621), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n457), .A2(new_n470), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(new_n418), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(new_n473), .A3(new_n474), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT90), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n626), .A2(new_n629), .A3(new_n630), .A4(new_n472), .ZN(new_n631));
  OAI21_X1  g430(.A(KEYINPUT37), .B1(new_n555), .B2(new_n559), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n610), .B1(new_n621), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n619), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n412), .A2(new_n410), .A3(new_n409), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n396), .A2(new_n406), .A3(G22gat), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n636), .B1(new_n637), .B2(new_n397), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n450), .B1(new_n440), .B2(new_n447), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT39), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n463), .A2(new_n436), .A3(new_n450), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT88), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n418), .B1(new_n639), .B2(new_n640), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT40), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n645), .A2(KEYINPUT40), .A3(new_n646), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n649), .A2(new_n628), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n638), .B1(new_n565), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n635), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n600), .A2(new_n602), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n638), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g455(.A(KEYINPUT35), .B1(new_n566), .B2(new_n656), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n562), .A2(new_n564), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n591), .A2(new_n594), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT35), .ZN(new_n662));
  NAND4_X1  g461(.A1(new_n661), .A2(new_n662), .A3(new_n609), .A4(new_n638), .ZN(new_n663));
  AOI22_X1  g462(.A1(new_n607), .A2(new_n654), .B1(new_n657), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT93), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n241), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n239), .A2(KEYINPUT93), .ZN(new_n667));
  OAI211_X1 g466(.A(new_n666), .B(new_n667), .C1(new_n287), .C2(new_n289), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n241), .A2(new_n242), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n239), .A2(KEYINPUT94), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n286), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(G229gat), .A2(G233gat), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n668), .A2(new_n671), .A3(KEYINPUT18), .A4(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n672), .B(KEYINPUT13), .Z(new_n674));
  INV_X1    g473(.A(new_n286), .ZN(new_n675));
  AND3_X1   g474(.A1(new_n243), .A2(new_n240), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n675), .B1(new_n243), .B2(new_n240), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n674), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n673), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT18), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT95), .ZN(new_n683));
  XNOR2_X1  g482(.A(G113gat), .B(G141gat), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G197gat), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT11), .B(G169gat), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(KEYINPUT91), .B(KEYINPUT12), .ZN(new_n688));
  XOR2_X1   g487(.A(new_n687), .B(new_n688), .Z(new_n689));
  OAI211_X1 g488(.A(new_n679), .B(new_n682), .C1(new_n683), .C2(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n673), .A2(new_n678), .A3(new_n683), .ZN(new_n691));
  INV_X1    g490(.A(new_n689), .ZN(new_n692));
  AND2_X1   g491(.A1(new_n680), .A2(new_n681), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n673), .A2(new_n678), .ZN(new_n694));
  OAI211_X1 g493(.A(new_n691), .B(new_n692), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  AND2_X1   g494(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n664), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT96), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n566), .A2(new_n413), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n604), .A2(new_n606), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g501(.A1(new_n626), .A2(new_n629), .A3(new_n472), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n633), .B1(new_n703), .B2(KEYINPUT90), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n652), .B1(new_n704), .B2(new_n631), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n638), .A2(new_n655), .ZN(new_n706));
  INV_X1    g505(.A(new_n608), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n628), .A2(KEYINPUT83), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n471), .A2(new_n475), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n658), .B1(new_n710), .B2(new_n472), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n662), .B1(new_n706), .B2(new_n711), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n609), .A2(new_n565), .A3(new_n659), .ZN(new_n713));
  NOR3_X1   g512(.A1(new_n713), .A2(new_n413), .A3(KEYINPUT35), .ZN(new_n714));
  OAI22_X1  g513(.A1(new_n702), .A2(new_n705), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n690), .A2(new_n695), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(KEYINPUT96), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n341), .B1(new_n699), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(new_n478), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(new_n232), .ZN(G1324gat));
  NOR2_X1   g520(.A1(new_n719), .A2(new_n565), .ZN(new_n722));
  XOR2_X1   g521(.A(KEYINPUT16), .B(G8gat), .Z(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(new_n238), .B2(new_n722), .ZN(new_n725));
  MUX2_X1   g524(.A(new_n724), .B(new_n725), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g525(.A(G15gat), .B1(new_n719), .B2(new_n701), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n660), .A2(G15gat), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n727), .B1(new_n719), .B2(new_n728), .ZN(G1326gat));
  OR3_X1    g528(.A1(new_n719), .A2(KEYINPUT107), .A3(new_n638), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT107), .B1(new_n719), .B2(new_n638), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT43), .B(G22gat), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(G1327gat));
  NOR2_X1   g533(.A1(new_n252), .A2(new_n340), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n735), .A2(new_n312), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n697), .A2(new_n698), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n717), .A2(KEYINPUT96), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n478), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n739), .A2(new_n278), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n741), .A2(KEYINPUT45), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n741), .A2(KEYINPUT45), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n664), .B2(new_n313), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n715), .A2(KEYINPUT44), .A3(new_n312), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n252), .A2(new_n696), .A3(new_n340), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G29gat), .B1(new_n749), .B2(new_n478), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n742), .B1(new_n743), .B2(new_n750), .ZN(G1328gat));
  NAND3_X1  g550(.A1(new_n739), .A2(new_n274), .A3(new_n658), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n752), .A2(KEYINPUT46), .ZN(new_n753));
  OAI21_X1  g552(.A(G36gat), .B1(new_n749), .B2(new_n565), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(KEYINPUT46), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(G1329gat));
  AOI21_X1  g555(.A(new_n605), .B1(new_n603), .B2(KEYINPUT36), .ZN(new_n757));
  AND4_X1   g556(.A1(G43gat), .A2(new_n747), .A3(new_n757), .A4(new_n748), .ZN(new_n758));
  AOI21_X1  g557(.A(G43gat), .B1(new_n739), .B2(new_n659), .ZN(new_n759));
  XNOR2_X1  g558(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n760));
  NOR4_X1   g559(.A1(new_n758), .A2(new_n759), .A3(KEYINPUT109), .A4(new_n760), .ZN(new_n761));
  NOR3_X1   g560(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT47), .B1(new_n758), .B2(new_n759), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n761), .B1(new_n764), .B2(new_n765), .ZN(G1330gat));
  INV_X1    g565(.A(G50gat), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n739), .A2(KEYINPUT110), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n413), .B1(new_n739), .B2(KEYINPUT110), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n767), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n413), .A2(G50gat), .ZN(new_n771));
  OR2_X1    g570(.A1(new_n749), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(KEYINPUT48), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n770), .A2(new_n775), .A3(new_n772), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n774), .A2(new_n776), .ZN(G1331gat));
  NOR2_X1   g576(.A1(new_n314), .A2(new_n716), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n340), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT111), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(new_n664), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(new_n740), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(G57gat), .ZN(G1332gat));
  INV_X1    g582(.A(new_n781), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n565), .ZN(new_n785));
  NOR2_X1   g584(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n786));
  AND2_X1   g585(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n788), .B1(new_n785), .B2(new_n786), .ZN(G1333gat));
  OAI21_X1  g588(.A(G71gat), .B1(new_n784), .B2(new_n701), .ZN(new_n790));
  INV_X1    g589(.A(G71gat), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n781), .A2(new_n791), .A3(new_n659), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT50), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n793), .B(new_n794), .ZN(G1334gat));
  NAND2_X1  g594(.A1(new_n781), .A2(new_n413), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G78gat), .ZN(G1335gat));
  INV_X1    g596(.A(new_n340), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n252), .A2(new_n716), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n745), .A2(new_n746), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(KEYINPUT112), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT112), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n745), .A2(new_n746), .A3(new_n802), .A4(new_n799), .ZN(new_n803));
  AND3_X1   g602(.A1(new_n801), .A2(new_n740), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g603(.A1(new_n664), .A2(new_n313), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n252), .A2(new_n716), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT51), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n805), .A2(KEYINPUT51), .A3(new_n806), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(new_n340), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n740), .A2(new_n254), .ZN(new_n813));
  OAI22_X1  g612(.A1(new_n804), .A2(new_n254), .B1(new_n812), .B2(new_n813), .ZN(G1336gat));
  NOR3_X1   g613(.A1(new_n798), .A2(G92gat), .A3(new_n565), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT113), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n811), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n253), .A2(new_n255), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n820), .B1(new_n800), .B2(new_n565), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n817), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n801), .A2(new_n658), .A3(new_n803), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n820), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n809), .A2(KEYINPUT114), .A3(new_n810), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT114), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n807), .A2(new_n827), .A3(new_n808), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n816), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n823), .B1(new_n830), .B2(KEYINPUT52), .ZN(new_n831));
  AOI211_X1 g630(.A(KEYINPUT115), .B(new_n818), .C1(new_n825), .C2(new_n829), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n822), .B1(new_n831), .B2(new_n832), .ZN(G1337gat));
  NAND3_X1  g632(.A1(new_n801), .A2(new_n757), .A3(new_n803), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT116), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n257), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n659), .A2(new_n257), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n812), .B2(new_n838), .ZN(G1338gat));
  NOR3_X1   g638(.A1(new_n798), .A2(new_n638), .A3(G106gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n811), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n842));
  OAI21_X1  g641(.A(G106gat), .B1(new_n800), .B2(new_n638), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n801), .A2(new_n413), .A3(new_n803), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT117), .ZN(new_n846));
  AND3_X1   g645(.A1(new_n845), .A2(new_n846), .A3(G106gat), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n845), .B2(G106gat), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n826), .A2(new_n828), .A3(new_n840), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n844), .B1(new_n850), .B2(new_n842), .ZN(G1339gat));
  NAND3_X1  g650(.A1(new_n679), .A2(new_n682), .A3(new_n689), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n676), .A2(new_n677), .A3(new_n674), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n672), .B1(new_n668), .B2(new_n671), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n687), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n856), .B1(new_n309), .B2(new_n311), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n334), .B1(new_n338), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n858), .B1(new_n323), .B2(new_n325), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n326), .A2(new_n861), .A3(new_n328), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT118), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n326), .A2(new_n861), .A3(KEYINPUT118), .A4(new_n328), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI22_X1  g665(.A1(new_n866), .A2(KEYINPUT55), .B1(new_n329), .B2(new_n336), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n857), .B(new_n867), .C1(KEYINPUT55), .C2(new_n866), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n798), .A2(new_n856), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n864), .A2(new_n865), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(new_n859), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT55), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n696), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n869), .B1(new_n873), .B2(new_n867), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n868), .B1(new_n874), .B2(new_n312), .ZN(new_n875));
  INV_X1    g674(.A(new_n252), .ZN(new_n876));
  AOI22_X1  g675(.A1(new_n875), .A2(new_n876), .B1(new_n798), .B2(new_n778), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n877), .A2(new_n478), .A3(new_n413), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n661), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n879), .A2(new_n422), .A3(new_n696), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n878), .A2(new_n565), .A3(new_n655), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n716), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n880), .B1(new_n882), .B2(new_n422), .ZN(G1340gat));
  NOR3_X1   g682(.A1(new_n879), .A2(new_n420), .A3(new_n798), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n340), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n885), .B2(new_n420), .ZN(G1341gat));
  NAND3_X1  g685(.A1(new_n881), .A2(new_n427), .A3(new_n252), .ZN(new_n887));
  OAI21_X1  g686(.A(G127gat), .B1(new_n879), .B2(new_n876), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(G1342gat));
  NAND2_X1  g688(.A1(new_n312), .A2(new_n565), .ZN(new_n890));
  XOR2_X1   g689(.A(new_n890), .B(KEYINPUT119), .Z(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n878), .A2(new_n425), .A3(new_n655), .A4(new_n892), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n893), .A2(KEYINPUT56), .ZN(new_n894));
  OAI21_X1  g693(.A(G134gat), .B1(new_n879), .B2(new_n313), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n893), .A2(KEYINPUT56), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(G1343gat));
  NOR2_X1   g696(.A1(new_n757), .A2(new_n478), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(new_n565), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n899), .B(KEYINPUT120), .Z(new_n900));
  INV_X1    g699(.A(KEYINPUT57), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n638), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n904), .B1(new_n874), .B2(new_n312), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n337), .B1(new_n871), .B2(new_n872), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n716), .B1(new_n866), .B2(KEYINPUT55), .ZN(new_n907));
  OAI22_X1  g706(.A1(new_n906), .A2(new_n907), .B1(new_n798), .B2(new_n856), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(KEYINPUT121), .A3(new_n313), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n905), .A2(new_n868), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n876), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n778), .A2(new_n798), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n903), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n875), .A2(new_n876), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n912), .ZN(new_n915));
  AOI21_X1  g714(.A(KEYINPUT57), .B1(new_n915), .B2(new_n413), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n716), .B(new_n900), .C1(new_n913), .C2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(KEYINPUT122), .B1(new_n917), .B2(G141gat), .ZN(new_n918));
  NAND4_X1  g717(.A1(new_n915), .A2(new_n413), .A3(new_n565), .A4(new_n898), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n919), .A2(G141gat), .A3(new_n696), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(new_n917), .B2(G141gat), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n918), .A2(new_n921), .A3(KEYINPUT58), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT58), .ZN(new_n923));
  AOI221_X4 g722(.A(new_n920), .B1(KEYINPUT122), .B2(new_n923), .C1(new_n917), .C2(G141gat), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n922), .A2(new_n924), .ZN(G1344gat));
  OAI21_X1  g724(.A(new_n901), .B1(new_n877), .B2(new_n638), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n915), .A2(new_n902), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n928), .A2(new_n340), .A3(new_n900), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n929), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n930));
  OAI21_X1  g729(.A(KEYINPUT59), .B1(new_n919), .B2(new_n798), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n931), .A2(new_n348), .A3(new_n350), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n913), .A2(new_n916), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT59), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n900), .A2(new_n934), .A3(new_n340), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n930), .B(new_n932), .C1(new_n933), .C2(new_n935), .ZN(G1345gat));
  OAI21_X1  g735(.A(new_n900), .B1(new_n913), .B2(new_n916), .ZN(new_n937));
  OAI21_X1  g736(.A(G155gat), .B1(new_n937), .B2(new_n876), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n252), .A2(new_n247), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n919), .B2(new_n939), .ZN(G1346gat));
  OAI21_X1  g739(.A(G162gat), .B1(new_n937), .B2(new_n313), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n915), .A2(new_n413), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n892), .A2(new_n361), .A3(new_n898), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(G1347gat));
  NOR2_X1   g743(.A1(new_n877), .A2(new_n413), .ZN(new_n945));
  NOR3_X1   g744(.A1(new_n740), .A2(new_n565), .A3(new_n660), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n947), .A2(new_n487), .A3(new_n696), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n656), .A2(new_n565), .ZN(new_n949));
  XNOR2_X1  g748(.A(new_n949), .B(KEYINPUT123), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n877), .A2(new_n740), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(G169gat), .B1(new_n951), .B2(new_n716), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n948), .A2(new_n952), .ZN(G1348gat));
  OAI21_X1  g752(.A(G176gat), .B1(new_n947), .B2(new_n798), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n951), .A2(new_n488), .A3(new_n340), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1349gat));
  OAI21_X1  g755(.A(G183gat), .B1(new_n947), .B2(new_n876), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n951), .A2(new_n530), .A3(new_n252), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT60), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n960), .A2(KEYINPUT124), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n959), .B(new_n961), .ZN(G1350gat));
  INV_X1    g761(.A(G190gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n951), .A2(new_n963), .A3(new_n312), .ZN(new_n964));
  OAI21_X1  g763(.A(G190gat), .B1(new_n947), .B2(new_n313), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n965), .A2(KEYINPUT61), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n965), .A2(KEYINPUT61), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(G1351gat));
  NAND3_X1  g767(.A1(new_n701), .A2(new_n413), .A3(new_n658), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n877), .A2(new_n740), .A3(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(G197gat), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n970), .A2(new_n971), .A3(new_n716), .ZN(new_n972));
  XOR2_X1   g771(.A(new_n972), .B(KEYINPUT125), .Z(new_n973));
  NOR2_X1   g772(.A1(new_n740), .A2(new_n565), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n701), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n975), .B1(new_n926), .B2(new_n927), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(G197gat), .B1(new_n977), .B2(new_n696), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n973), .A2(new_n978), .ZN(G1352gat));
  OAI21_X1  g778(.A(G204gat), .B1(new_n977), .B2(new_n798), .ZN(new_n980));
  INV_X1    g779(.A(G204gat), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n970), .A2(new_n981), .A3(new_n340), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT62), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n983), .A2(KEYINPUT126), .ZN(new_n984));
  AND2_X1   g783(.A1(new_n983), .A2(KEYINPUT126), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI211_X1 g785(.A(new_n980), .B(new_n986), .C1(new_n984), .C2(new_n982), .ZN(G1353gat));
  INV_X1    g786(.A(KEYINPUT63), .ZN(new_n988));
  INV_X1    g787(.A(new_n975), .ZN(new_n989));
  NOR2_X1   g788(.A1(new_n877), .A2(new_n903), .ZN(new_n990));
  OAI211_X1 g789(.A(new_n252), .B(new_n989), .C1(new_n916), .C2(new_n990), .ZN(new_n991));
  OAI21_X1  g790(.A(G211gat), .B1(new_n991), .B2(KEYINPUT127), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n993));
  AOI21_X1  g792(.A(new_n993), .B1(new_n976), .B2(new_n252), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n988), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n991), .A2(KEYINPUT127), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n976), .A2(new_n993), .A3(new_n252), .ZN(new_n997));
  NAND4_X1  g796(.A1(new_n996), .A2(KEYINPUT63), .A3(new_n997), .A4(G211gat), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n970), .A2(new_n371), .A3(new_n252), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(G1354gat));
  OAI21_X1  g800(.A(G218gat), .B1(new_n977), .B2(new_n313), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n970), .A2(new_n372), .A3(new_n312), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(G1355gat));
endmodule


