

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U546 ( .A(n645), .B(n590), .ZN(n630) );
  NOR2_X2 U547 ( .A1(G2104), .A2(n522), .ZN(n882) );
  INV_X1 U548 ( .A(G2105), .ZN(n522) );
  NOR2_X2 U549 ( .A1(n525), .A2(n524), .ZN(n584) );
  NOR2_X1 U550 ( .A1(G2105), .A2(G2104), .ZN(n517) );
  NOR2_X1 U551 ( .A1(n663), .A2(n847), .ZN(n605) );
  INV_X1 U552 ( .A(KEYINPUT26), .ZN(n604) );
  NOR2_X1 U553 ( .A1(G1384), .A2(G164), .ZN(n588) );
  AND2_X1 U554 ( .A1(n618), .A2(n617), .ZN(n635) );
  XNOR2_X1 U555 ( .A(n586), .B(n585), .ZN(n729) );
  AND2_X1 U556 ( .A1(n963), .A2(n512), .ZN(n682) );
  BUF_X1 U557 ( .A(n526), .Z(n877) );
  AND2_X1 U558 ( .A1(n526), .A2(G137), .ZN(n519) );
  NOR2_X1 U559 ( .A1(n533), .A2(n532), .ZN(G164) );
  BUF_X1 U560 ( .A(n584), .Z(G160) );
  AND2_X1 U561 ( .A1(n688), .A2(n687), .ZN(n510) );
  XOR2_X1 U562 ( .A(KEYINPUT40), .B(KEYINPUT104), .Z(n511) );
  OR2_X1 U563 ( .A1(G1971), .A2(G303), .ZN(n512) );
  INV_X1 U564 ( .A(KEYINPUT95), .ZN(n591) );
  XNOR2_X1 U565 ( .A(n592), .B(n591), .ZN(n595) );
  INV_X1 U566 ( .A(n964), .ZN(n615) );
  AND2_X1 U567 ( .A1(n616), .A2(n615), .ZN(n617) );
  AND2_X1 U568 ( .A1(n637), .A2(n636), .ZN(n638) );
  INV_X1 U569 ( .A(KEYINPUT98), .ZN(n650) );
  INV_X1 U570 ( .A(KEYINPUT92), .ZN(n587) );
  INV_X1 U571 ( .A(n645), .ZN(n663) );
  AND2_X1 U572 ( .A1(n670), .A2(n669), .ZN(n672) );
  INV_X1 U573 ( .A(n744), .ZN(n687) );
  INV_X1 U574 ( .A(KEYINPUT17), .ZN(n516) );
  XNOR2_X1 U575 ( .A(n517), .B(n516), .ZN(n526) );
  NOR2_X1 U576 ( .A1(G543), .A2(G651), .ZN(n795) );
  NOR2_X1 U577 ( .A1(n567), .A2(G651), .ZN(n799) );
  AND2_X4 U578 ( .A1(n522), .A2(G2104), .ZN(n876) );
  NAND2_X1 U579 ( .A1(G101), .A2(n876), .ZN(n513) );
  XOR2_X1 U580 ( .A(n513), .B(KEYINPUT23), .Z(n515) );
  AND2_X1 U581 ( .A1(G2105), .A2(G2104), .ZN(n881) );
  NAND2_X1 U582 ( .A1(n881), .A2(G113), .ZN(n514) );
  AND2_X1 U583 ( .A1(n515), .A2(n514), .ZN(n521) );
  INV_X1 U584 ( .A(KEYINPUT66), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n519), .B(n518), .ZN(n520) );
  NAND2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n525) );
  NAND2_X1 U587 ( .A1(G125), .A2(n882), .ZN(n523) );
  XNOR2_X1 U588 ( .A(KEYINPUT65), .B(n523), .ZN(n524) );
  NAND2_X1 U589 ( .A1(G102), .A2(n876), .ZN(n528) );
  NAND2_X1 U590 ( .A1(G138), .A2(n526), .ZN(n527) );
  NAND2_X1 U591 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U592 ( .A(KEYINPUT84), .B(n529), .ZN(n533) );
  NAND2_X1 U593 ( .A1(G114), .A2(n881), .ZN(n531) );
  NAND2_X1 U594 ( .A1(G126), .A2(n882), .ZN(n530) );
  NAND2_X1 U595 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U596 ( .A1(n795), .A2(G90), .ZN(n534) );
  XNOR2_X1 U597 ( .A(n534), .B(KEYINPUT68), .ZN(n536) );
  XOR2_X1 U598 ( .A(KEYINPUT0), .B(G543), .Z(n567) );
  XNOR2_X1 U599 ( .A(KEYINPUT67), .B(G651), .ZN(n538) );
  NOR2_X1 U600 ( .A1(n567), .A2(n538), .ZN(n800) );
  NAND2_X1 U601 ( .A1(G77), .A2(n800), .ZN(n535) );
  NAND2_X1 U602 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U603 ( .A(KEYINPUT9), .B(n537), .ZN(n543) );
  NOR2_X1 U604 ( .A1(G543), .A2(n538), .ZN(n539) );
  XOR2_X1 U605 ( .A(KEYINPUT1), .B(n539), .Z(n796) );
  NAND2_X1 U606 ( .A1(n796), .A2(G64), .ZN(n541) );
  NAND2_X1 U607 ( .A1(n799), .A2(G52), .ZN(n540) );
  AND2_X1 U608 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U609 ( .A1(n543), .A2(n542), .ZN(G301) );
  NAND2_X1 U610 ( .A1(n799), .A2(G51), .ZN(n545) );
  NAND2_X1 U611 ( .A1(G63), .A2(n796), .ZN(n544) );
  NAND2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(KEYINPUT6), .B(n546), .ZN(n552) );
  NAND2_X1 U614 ( .A1(n795), .A2(G89), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n547), .B(KEYINPUT4), .ZN(n549) );
  NAND2_X1 U616 ( .A1(G76), .A2(n800), .ZN(n548) );
  NAND2_X1 U617 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U618 ( .A(n550), .B(KEYINPUT5), .Z(n551) );
  NOR2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U620 ( .A(KEYINPUT7), .B(n553), .Z(n554) );
  XOR2_X1 U621 ( .A(KEYINPUT73), .B(n554), .Z(G168) );
  XOR2_X1 U622 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U623 ( .A1(G88), .A2(n795), .ZN(n555) );
  XNOR2_X1 U624 ( .A(n555), .B(KEYINPUT82), .ZN(n562) );
  NAND2_X1 U625 ( .A1(G62), .A2(n796), .ZN(n557) );
  NAND2_X1 U626 ( .A1(G75), .A2(n800), .ZN(n556) );
  NAND2_X1 U627 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U628 ( .A1(G50), .A2(n799), .ZN(n558) );
  XNOR2_X1 U629 ( .A(KEYINPUT81), .B(n558), .ZN(n559) );
  NOR2_X1 U630 ( .A1(n560), .A2(n559), .ZN(n561) );
  NAND2_X1 U631 ( .A1(n562), .A2(n561), .ZN(G303) );
  NAND2_X1 U632 ( .A1(G49), .A2(n799), .ZN(n564) );
  NAND2_X1 U633 ( .A1(G74), .A2(G651), .ZN(n563) );
  NAND2_X1 U634 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U635 ( .A1(n796), .A2(n565), .ZN(n566) );
  XOR2_X1 U636 ( .A(KEYINPUT79), .B(n566), .Z(n569) );
  NAND2_X1 U637 ( .A1(n567), .A2(G87), .ZN(n568) );
  NAND2_X1 U638 ( .A1(n569), .A2(n568), .ZN(G288) );
  NAND2_X1 U639 ( .A1(G86), .A2(n795), .ZN(n570) );
  XNOR2_X1 U640 ( .A(n570), .B(KEYINPUT80), .ZN(n577) );
  NAND2_X1 U641 ( .A1(n799), .A2(G48), .ZN(n572) );
  NAND2_X1 U642 ( .A1(G61), .A2(n796), .ZN(n571) );
  NAND2_X1 U643 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U644 ( .A1(n800), .A2(G73), .ZN(n573) );
  XOR2_X1 U645 ( .A(KEYINPUT2), .B(n573), .Z(n574) );
  NOR2_X1 U646 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U647 ( .A1(n577), .A2(n576), .ZN(G305) );
  NAND2_X1 U648 ( .A1(n795), .A2(G85), .ZN(n579) );
  NAND2_X1 U649 ( .A1(G60), .A2(n796), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n579), .A2(n578), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n799), .A2(G47), .ZN(n581) );
  NAND2_X1 U652 ( .A1(G72), .A2(n800), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n581), .A2(n580), .ZN(n582) );
  OR2_X1 U654 ( .A1(n583), .A2(n582), .ZN(G290) );
  NAND2_X1 U655 ( .A1(G40), .A2(n584), .ZN(n586) );
  INV_X1 U656 ( .A(KEYINPUT85), .ZN(n585) );
  XNOR2_X1 U657 ( .A(n729), .B(n587), .ZN(n589) );
  XNOR2_X1 U658 ( .A(n588), .B(KEYINPUT64), .ZN(n730) );
  AND2_X2 U659 ( .A1(n589), .A2(n730), .ZN(n645) );
  INV_X1 U660 ( .A(KEYINPUT93), .ZN(n590) );
  NAND2_X1 U661 ( .A1(G2067), .A2(n630), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G1348), .A2(n663), .ZN(n593) );
  XNOR2_X1 U663 ( .A(KEYINPUT94), .B(n593), .ZN(n594) );
  NAND2_X1 U664 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U665 ( .A(n596), .B(KEYINPUT96), .ZN(n620) );
  NAND2_X1 U666 ( .A1(n795), .A2(G92), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G66), .A2(n796), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U669 ( .A1(n799), .A2(G54), .ZN(n600) );
  NAND2_X1 U670 ( .A1(G79), .A2(n800), .ZN(n599) );
  NAND2_X1 U671 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U672 ( .A1(n602), .A2(n601), .ZN(n603) );
  XOR2_X1 U673 ( .A(KEYINPUT15), .B(n603), .Z(n971) );
  INV_X1 U674 ( .A(G1996), .ZN(n847) );
  XNOR2_X1 U675 ( .A(n605), .B(n604), .ZN(n618) );
  NAND2_X1 U676 ( .A1(n663), .A2(G1341), .ZN(n616) );
  NAND2_X1 U677 ( .A1(n796), .A2(G56), .ZN(n606) );
  XOR2_X1 U678 ( .A(KEYINPUT14), .B(n606), .Z(n612) );
  NAND2_X1 U679 ( .A1(n795), .A2(G81), .ZN(n607) );
  XNOR2_X1 U680 ( .A(n607), .B(KEYINPUT12), .ZN(n609) );
  NAND2_X1 U681 ( .A1(G68), .A2(n800), .ZN(n608) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n610) );
  XOR2_X1 U683 ( .A(KEYINPUT13), .B(n610), .Z(n611) );
  NOR2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n799), .A2(G43), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n964) );
  NOR2_X1 U687 ( .A1(n971), .A2(n635), .ZN(n619) );
  NOR2_X1 U688 ( .A1(n620), .A2(n619), .ZN(n634) );
  NAND2_X1 U689 ( .A1(n800), .A2(G78), .ZN(n627) );
  NAND2_X1 U690 ( .A1(n795), .A2(G91), .ZN(n622) );
  NAND2_X1 U691 ( .A1(G65), .A2(n796), .ZN(n621) );
  NAND2_X1 U692 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U693 ( .A1(G53), .A2(n799), .ZN(n623) );
  XNOR2_X1 U694 ( .A(KEYINPUT69), .B(n623), .ZN(n624) );
  NOR2_X1 U695 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U697 ( .A(n628), .B(KEYINPUT70), .ZN(n972) );
  NAND2_X1 U698 ( .A1(n630), .A2(G2072), .ZN(n629) );
  XOR2_X1 U699 ( .A(KEYINPUT27), .B(n629), .Z(n632) );
  INV_X1 U700 ( .A(n630), .ZN(n644) );
  NAND2_X1 U701 ( .A1(G1956), .A2(n644), .ZN(n631) );
  NAND2_X1 U702 ( .A1(n632), .A2(n631), .ZN(n639) );
  NOR2_X1 U703 ( .A1(n972), .A2(n639), .ZN(n633) );
  NOR2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U705 ( .A1(n971), .A2(n635), .ZN(n636) );
  XNOR2_X1 U706 ( .A(n638), .B(KEYINPUT97), .ZN(n642) );
  NAND2_X1 U707 ( .A1(n972), .A2(n639), .ZN(n640) );
  XNOR2_X1 U708 ( .A(KEYINPUT28), .B(n640), .ZN(n641) );
  NAND2_X1 U709 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X1 U710 ( .A(n643), .B(KEYINPUT29), .ZN(n649) );
  XOR2_X1 U711 ( .A(KEYINPUT25), .B(G2078), .Z(n943) );
  NOR2_X1 U712 ( .A1(n943), .A2(n644), .ZN(n647) );
  NOR2_X1 U713 ( .A1(n645), .A2(G1961), .ZN(n646) );
  NOR2_X1 U714 ( .A1(n647), .A2(n646), .ZN(n652) );
  NOR2_X1 U715 ( .A1(G301), .A2(n652), .ZN(n648) );
  NOR2_X2 U716 ( .A1(n649), .A2(n648), .ZN(n651) );
  XNOR2_X1 U717 ( .A(n651), .B(n650), .ZN(n661) );
  AND2_X1 U718 ( .A1(G301), .A2(n652), .ZN(n657) );
  NAND2_X1 U719 ( .A1(G8), .A2(n663), .ZN(n744) );
  NOR2_X1 U720 ( .A1(G1966), .A2(n744), .ZN(n676) );
  NOR2_X1 U721 ( .A1(G2084), .A2(n663), .ZN(n673) );
  NOR2_X1 U722 ( .A1(n676), .A2(n673), .ZN(n653) );
  NAND2_X1 U723 ( .A1(G8), .A2(n653), .ZN(n654) );
  XNOR2_X1 U724 ( .A(KEYINPUT30), .B(n654), .ZN(n655) );
  NOR2_X1 U725 ( .A1(G168), .A2(n655), .ZN(n656) );
  NOR2_X1 U726 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U727 ( .A(KEYINPUT31), .B(n658), .ZN(n659) );
  XNOR2_X1 U728 ( .A(n659), .B(KEYINPUT99), .ZN(n660) );
  NAND2_X1 U729 ( .A1(n661), .A2(n660), .ZN(n674) );
  XNOR2_X1 U730 ( .A(n674), .B(KEYINPUT100), .ZN(n662) );
  NAND2_X1 U731 ( .A1(n662), .A2(G286), .ZN(n670) );
  INV_X1 U732 ( .A(G8), .ZN(n668) );
  NOR2_X1 U733 ( .A1(G1971), .A2(n744), .ZN(n665) );
  NOR2_X1 U734 ( .A1(G2090), .A2(n663), .ZN(n664) );
  NOR2_X1 U735 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U736 ( .A1(n666), .A2(G303), .ZN(n667) );
  OR2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U738 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n671) );
  XNOR2_X1 U739 ( .A(n672), .B(n671), .ZN(n680) );
  NAND2_X1 U740 ( .A1(G8), .A2(n673), .ZN(n678) );
  XOR2_X1 U741 ( .A(KEYINPUT100), .B(n674), .Z(n675) );
  NOR2_X1 U742 ( .A1(n676), .A2(n675), .ZN(n677) );
  NAND2_X1 U743 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U744 ( .A1(n680), .A2(n679), .ZN(n734) );
  NOR2_X1 U745 ( .A1(G288), .A2(G1976), .ZN(n681) );
  XOR2_X1 U746 ( .A(n681), .B(KEYINPUT102), .Z(n963) );
  NAND2_X1 U747 ( .A1(n734), .A2(n682), .ZN(n689) );
  NAND2_X1 U748 ( .A1(G1976), .A2(G288), .ZN(n969) );
  INV_X1 U749 ( .A(KEYINPUT33), .ZN(n739) );
  OR2_X1 U750 ( .A1(n744), .A2(n963), .ZN(n683) );
  NOR2_X1 U751 ( .A1(n739), .A2(n683), .ZN(n684) );
  XNOR2_X1 U752 ( .A(n684), .B(KEYINPUT103), .ZN(n738) );
  AND2_X1 U753 ( .A1(n969), .A2(n738), .ZN(n686) );
  XNOR2_X1 U754 ( .A(G1981), .B(G305), .ZN(n980) );
  INV_X1 U755 ( .A(n980), .ZN(n685) );
  AND2_X1 U756 ( .A1(n686), .A2(n685), .ZN(n688) );
  NAND2_X1 U757 ( .A1(n689), .A2(n510), .ZN(n750) );
  NOR2_X1 U758 ( .A1(G2090), .A2(G303), .ZN(n690) );
  NAND2_X1 U759 ( .A1(G8), .A2(n690), .ZN(n732) );
  NAND2_X1 U760 ( .A1(G129), .A2(n882), .ZN(n692) );
  NAND2_X1 U761 ( .A1(G141), .A2(n877), .ZN(n691) );
  NAND2_X1 U762 ( .A1(n692), .A2(n691), .ZN(n695) );
  NAND2_X1 U763 ( .A1(n876), .A2(G105), .ZN(n693) );
  XOR2_X1 U764 ( .A(KEYINPUT38), .B(n693), .Z(n694) );
  NOR2_X1 U765 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U766 ( .A1(n881), .A2(G117), .ZN(n696) );
  NAND2_X1 U767 ( .A1(n697), .A2(n696), .ZN(n895) );
  NOR2_X1 U768 ( .A1(G1996), .A2(n895), .ZN(n989) );
  NAND2_X1 U769 ( .A1(G119), .A2(n882), .ZN(n699) );
  NAND2_X1 U770 ( .A1(G95), .A2(n876), .ZN(n698) );
  NAND2_X1 U771 ( .A1(n699), .A2(n698), .ZN(n704) );
  NAND2_X1 U772 ( .A1(n881), .A2(G107), .ZN(n700) );
  XNOR2_X1 U773 ( .A(n700), .B(KEYINPUT88), .ZN(n702) );
  NAND2_X1 U774 ( .A1(G131), .A2(n877), .ZN(n701) );
  NAND2_X1 U775 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U776 ( .A1(n704), .A2(n703), .ZN(n705) );
  XNOR2_X1 U777 ( .A(n705), .B(KEYINPUT89), .ZN(n890) );
  NAND2_X1 U778 ( .A1(G1991), .A2(n890), .ZN(n706) );
  XNOR2_X1 U779 ( .A(KEYINPUT90), .B(n706), .ZN(n709) );
  NAND2_X1 U780 ( .A1(G1996), .A2(n895), .ZN(n707) );
  XOR2_X1 U781 ( .A(KEYINPUT91), .B(n707), .Z(n708) );
  NAND2_X1 U782 ( .A1(n709), .A2(n708), .ZN(n751) );
  NOR2_X1 U783 ( .A1(G1986), .A2(G290), .ZN(n710) );
  NOR2_X1 U784 ( .A1(G1991), .A2(n890), .ZN(n995) );
  NOR2_X1 U785 ( .A1(n710), .A2(n995), .ZN(n711) );
  NOR2_X1 U786 ( .A1(n751), .A2(n711), .ZN(n712) );
  NOR2_X1 U787 ( .A1(n989), .A2(n712), .ZN(n713) );
  XNOR2_X1 U788 ( .A(KEYINPUT39), .B(n713), .ZN(n726) );
  XNOR2_X1 U789 ( .A(G2067), .B(KEYINPUT37), .ZN(n714) );
  XNOR2_X1 U790 ( .A(n714), .B(KEYINPUT86), .ZN(n727) );
  NAND2_X1 U791 ( .A1(n876), .A2(G104), .ZN(n715) );
  XOR2_X1 U792 ( .A(KEYINPUT87), .B(n715), .Z(n717) );
  NAND2_X1 U793 ( .A1(n877), .A2(G140), .ZN(n716) );
  NAND2_X1 U794 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U795 ( .A(KEYINPUT34), .B(n718), .ZN(n723) );
  NAND2_X1 U796 ( .A1(G116), .A2(n881), .ZN(n720) );
  NAND2_X1 U797 ( .A1(G128), .A2(n882), .ZN(n719) );
  NAND2_X1 U798 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U799 ( .A(KEYINPUT35), .B(n721), .Z(n722) );
  NOR2_X1 U800 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U801 ( .A(KEYINPUT36), .B(n724), .ZN(n898) );
  NOR2_X1 U802 ( .A1(n727), .A2(n898), .ZN(n752) );
  INV_X1 U803 ( .A(n752), .ZN(n725) );
  NAND2_X1 U804 ( .A1(n726), .A2(n725), .ZN(n728) );
  NAND2_X1 U805 ( .A1(n727), .A2(n898), .ZN(n991) );
  NAND2_X1 U806 ( .A1(n728), .A2(n991), .ZN(n731) );
  NOR2_X1 U807 ( .A1(n730), .A2(n729), .ZN(n753) );
  NAND2_X1 U808 ( .A1(n731), .A2(n753), .ZN(n735) );
  AND2_X1 U809 ( .A1(n732), .A2(n735), .ZN(n733) );
  NAND2_X1 U810 ( .A1(n734), .A2(n733), .ZN(n737) );
  INV_X1 U811 ( .A(n735), .ZN(n756) );
  OR2_X1 U812 ( .A1(n756), .A2(n744), .ZN(n736) );
  NAND2_X1 U813 ( .A1(n737), .A2(n736), .ZN(n748) );
  INV_X1 U814 ( .A(n738), .ZN(n740) );
  OR2_X1 U815 ( .A1(n740), .A2(n739), .ZN(n741) );
  NOR2_X1 U816 ( .A1(n980), .A2(n741), .ZN(n746) );
  NOR2_X1 U817 ( .A1(G1981), .A2(G305), .ZN(n742) );
  XOR2_X1 U818 ( .A(n742), .B(KEYINPUT24), .Z(n743) );
  NOR2_X1 U819 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U820 ( .A1(n746), .A2(n745), .ZN(n747) );
  AND2_X1 U821 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U822 ( .A1(n750), .A2(n749), .ZN(n758) );
  XOR2_X1 U823 ( .A(G1986), .B(G290), .Z(n970) );
  NOR2_X1 U824 ( .A1(n752), .A2(n751), .ZN(n1001) );
  NAND2_X1 U825 ( .A1(n970), .A2(n1001), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n754), .A2(n753), .ZN(n755) );
  OR2_X1 U827 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U828 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U829 ( .A(n759), .B(n511), .ZN(G329) );
  XOR2_X1 U830 ( .A(G2435), .B(G2454), .Z(n761) );
  XNOR2_X1 U831 ( .A(KEYINPUT105), .B(G2438), .ZN(n760) );
  XNOR2_X1 U832 ( .A(n761), .B(n760), .ZN(n768) );
  XOR2_X1 U833 ( .A(G2446), .B(G2430), .Z(n763) );
  XNOR2_X1 U834 ( .A(G2451), .B(G2443), .ZN(n762) );
  XNOR2_X1 U835 ( .A(n763), .B(n762), .ZN(n764) );
  XOR2_X1 U836 ( .A(n764), .B(G2427), .Z(n766) );
  XNOR2_X1 U837 ( .A(G1341), .B(G1348), .ZN(n765) );
  XNOR2_X1 U838 ( .A(n766), .B(n765), .ZN(n767) );
  XNOR2_X1 U839 ( .A(n768), .B(n767), .ZN(n769) );
  AND2_X1 U840 ( .A1(n769), .A2(G14), .ZN(G401) );
  AND2_X1 U841 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U842 ( .A(G57), .ZN(G237) );
  INV_X1 U843 ( .A(G82), .ZN(G220) );
  NAND2_X1 U844 ( .A1(G7), .A2(G661), .ZN(n770) );
  XOR2_X1 U845 ( .A(n770), .B(KEYINPUT10), .Z(n915) );
  NAND2_X1 U846 ( .A1(n915), .A2(G567), .ZN(n771) );
  XOR2_X1 U847 ( .A(KEYINPUT11), .B(n771), .Z(G234) );
  INV_X1 U848 ( .A(G860), .ZN(n776) );
  OR2_X1 U849 ( .A1(n964), .A2(n776), .ZN(G153) );
  NAND2_X1 U850 ( .A1(G868), .A2(G301), .ZN(n773) );
  OR2_X1 U851 ( .A1(n971), .A2(G868), .ZN(n772) );
  NAND2_X1 U852 ( .A1(n773), .A2(n772), .ZN(G284) );
  XOR2_X1 U853 ( .A(n972), .B(KEYINPUT71), .Z(G299) );
  NOR2_X1 U854 ( .A1(G868), .A2(G299), .ZN(n775) );
  INV_X1 U855 ( .A(G868), .ZN(n815) );
  NOR2_X1 U856 ( .A1(G286), .A2(n815), .ZN(n774) );
  NOR2_X1 U857 ( .A1(n775), .A2(n774), .ZN(G297) );
  NAND2_X1 U858 ( .A1(n776), .A2(G559), .ZN(n777) );
  NAND2_X1 U859 ( .A1(n777), .A2(n971), .ZN(n778) );
  XNOR2_X1 U860 ( .A(n778), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U861 ( .A1(G868), .A2(n964), .ZN(n781) );
  NAND2_X1 U862 ( .A1(G868), .A2(n971), .ZN(n779) );
  NOR2_X1 U863 ( .A1(G559), .A2(n779), .ZN(n780) );
  NOR2_X1 U864 ( .A1(n781), .A2(n780), .ZN(G282) );
  NAND2_X1 U865 ( .A1(G111), .A2(n881), .ZN(n783) );
  NAND2_X1 U866 ( .A1(G135), .A2(n877), .ZN(n782) );
  NAND2_X1 U867 ( .A1(n783), .A2(n782), .ZN(n788) );
  XOR2_X1 U868 ( .A(KEYINPUT18), .B(KEYINPUT75), .Z(n785) );
  NAND2_X1 U869 ( .A1(G123), .A2(n882), .ZN(n784) );
  XNOR2_X1 U870 ( .A(n785), .B(n784), .ZN(n786) );
  XOR2_X1 U871 ( .A(KEYINPUT74), .B(n786), .Z(n787) );
  NOR2_X1 U872 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U873 ( .A1(n876), .A2(G99), .ZN(n789) );
  NAND2_X1 U874 ( .A1(n790), .A2(n789), .ZN(n993) );
  XNOR2_X1 U875 ( .A(n993), .B(G2096), .ZN(n792) );
  XNOR2_X1 U876 ( .A(G2100), .B(KEYINPUT76), .ZN(n791) );
  NOR2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n793) );
  XNOR2_X1 U878 ( .A(KEYINPUT77), .B(n793), .ZN(G156) );
  NAND2_X1 U879 ( .A1(G559), .A2(n971), .ZN(n794) );
  XNOR2_X1 U880 ( .A(n794), .B(n964), .ZN(n812) );
  NOR2_X1 U881 ( .A1(G860), .A2(n812), .ZN(n806) );
  NAND2_X1 U882 ( .A1(n795), .A2(G93), .ZN(n798) );
  NAND2_X1 U883 ( .A1(G67), .A2(n796), .ZN(n797) );
  NAND2_X1 U884 ( .A1(n798), .A2(n797), .ZN(n804) );
  NAND2_X1 U885 ( .A1(n799), .A2(G55), .ZN(n802) );
  NAND2_X1 U886 ( .A1(G80), .A2(n800), .ZN(n801) );
  NAND2_X1 U887 ( .A1(n802), .A2(n801), .ZN(n803) );
  OR2_X1 U888 ( .A1(n804), .A2(n803), .ZN(n814) );
  XOR2_X1 U889 ( .A(n814), .B(KEYINPUT78), .Z(n805) );
  XNOR2_X1 U890 ( .A(n806), .B(n805), .ZN(G145) );
  XOR2_X1 U891 ( .A(G303), .B(KEYINPUT19), .Z(n811) );
  XOR2_X1 U892 ( .A(n814), .B(G290), .Z(n809) );
  XOR2_X1 U893 ( .A(G299), .B(G305), .Z(n807) );
  XNOR2_X1 U894 ( .A(G288), .B(n807), .ZN(n808) );
  XNOR2_X1 U895 ( .A(n809), .B(n808), .ZN(n810) );
  XNOR2_X1 U896 ( .A(n811), .B(n810), .ZN(n901) );
  XNOR2_X1 U897 ( .A(n812), .B(n901), .ZN(n813) );
  NAND2_X1 U898 ( .A1(n813), .A2(G868), .ZN(n817) );
  NAND2_X1 U899 ( .A1(n815), .A2(n814), .ZN(n816) );
  NAND2_X1 U900 ( .A1(n817), .A2(n816), .ZN(G295) );
  XOR2_X1 U901 ( .A(KEYINPUT21), .B(KEYINPUT83), .Z(n821) );
  NAND2_X1 U902 ( .A1(G2084), .A2(G2078), .ZN(n818) );
  XOR2_X1 U903 ( .A(KEYINPUT20), .B(n818), .Z(n819) );
  NAND2_X1 U904 ( .A1(n819), .A2(G2090), .ZN(n820) );
  XNOR2_X1 U905 ( .A(n821), .B(n820), .ZN(n822) );
  NAND2_X1 U906 ( .A1(G2072), .A2(n822), .ZN(G158) );
  XNOR2_X1 U907 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U908 ( .A(KEYINPUT72), .B(G132), .Z(G219) );
  NOR2_X1 U909 ( .A1(G219), .A2(G220), .ZN(n823) );
  XOR2_X1 U910 ( .A(KEYINPUT22), .B(n823), .Z(n824) );
  NOR2_X1 U911 ( .A1(G218), .A2(n824), .ZN(n825) );
  NAND2_X1 U912 ( .A1(G96), .A2(n825), .ZN(n834) );
  NAND2_X1 U913 ( .A1(n834), .A2(G2106), .ZN(n829) );
  NAND2_X1 U914 ( .A1(G108), .A2(G120), .ZN(n826) );
  NOR2_X1 U915 ( .A1(G237), .A2(n826), .ZN(n827) );
  NAND2_X1 U916 ( .A1(G69), .A2(n827), .ZN(n835) );
  NAND2_X1 U917 ( .A1(n835), .A2(G567), .ZN(n828) );
  NAND2_X1 U918 ( .A1(n829), .A2(n828), .ZN(n914) );
  NAND2_X1 U919 ( .A1(G661), .A2(G483), .ZN(n830) );
  NOR2_X1 U920 ( .A1(n914), .A2(n830), .ZN(n833) );
  NAND2_X1 U921 ( .A1(n833), .A2(G36), .ZN(G176) );
  NAND2_X1 U922 ( .A1(G2106), .A2(n915), .ZN(G217) );
  AND2_X1 U923 ( .A1(G15), .A2(G2), .ZN(n831) );
  NAND2_X1 U924 ( .A1(G661), .A2(n831), .ZN(G259) );
  NAND2_X1 U925 ( .A1(G3), .A2(G1), .ZN(n832) );
  NAND2_X1 U926 ( .A1(n833), .A2(n832), .ZN(G188) );
  XOR2_X1 U927 ( .A(G120), .B(KEYINPUT106), .Z(G236) );
  INV_X1 U929 ( .A(G108), .ZN(G238) );
  INV_X1 U930 ( .A(G96), .ZN(G221) );
  NOR2_X1 U931 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U932 ( .A(G325), .ZN(G261) );
  XOR2_X1 U933 ( .A(KEYINPUT42), .B(G2090), .Z(n837) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2078), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U936 ( .A(n838), .B(G2100), .Z(n840) );
  XNOR2_X1 U937 ( .A(G2084), .B(G2072), .ZN(n839) );
  XNOR2_X1 U938 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U939 ( .A(G2096), .B(KEYINPUT43), .Z(n842) );
  XNOR2_X1 U940 ( .A(KEYINPUT107), .B(G2678), .ZN(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U942 ( .A(n844), .B(n843), .Z(G227) );
  XOR2_X1 U943 ( .A(G1976), .B(G1981), .Z(n846) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1971), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n857) );
  XOR2_X1 U946 ( .A(KEYINPUT41), .B(G2474), .Z(n849) );
  XOR2_X1 U947 ( .A(n847), .B(KEYINPUT108), .Z(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U949 ( .A(G1956), .B(G1961), .Z(n851) );
  XNOR2_X1 U950 ( .A(G1991), .B(G1986), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U952 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U953 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U955 ( .A(n857), .B(n856), .ZN(G229) );
  NAND2_X1 U956 ( .A1(G124), .A2(n882), .ZN(n858) );
  XNOR2_X1 U957 ( .A(n858), .B(KEYINPUT44), .ZN(n861) );
  NAND2_X1 U958 ( .A1(G100), .A2(n876), .ZN(n859) );
  XOR2_X1 U959 ( .A(KEYINPUT111), .B(n859), .Z(n860) );
  NAND2_X1 U960 ( .A1(n861), .A2(n860), .ZN(n865) );
  NAND2_X1 U961 ( .A1(G112), .A2(n881), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G136), .A2(n877), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n864) );
  NOR2_X1 U964 ( .A1(n865), .A2(n864), .ZN(G162) );
  NAND2_X1 U965 ( .A1(G130), .A2(n882), .ZN(n874) );
  XNOR2_X1 U966 ( .A(KEYINPUT113), .B(KEYINPUT45), .ZN(n869) );
  NAND2_X1 U967 ( .A1(G106), .A2(n876), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G142), .A2(n877), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n869), .B(n868), .ZN(n872) );
  NAND2_X1 U971 ( .A1(n881), .A2(G118), .ZN(n870) );
  XOR2_X1 U972 ( .A(KEYINPUT112), .B(n870), .Z(n871) );
  NOR2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n873) );
  NAND2_X1 U974 ( .A1(n874), .A2(n873), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n875), .B(KEYINPUT46), .ZN(n894) );
  NAND2_X1 U976 ( .A1(G103), .A2(n876), .ZN(n879) );
  NAND2_X1 U977 ( .A1(G139), .A2(n877), .ZN(n878) );
  NAND2_X1 U978 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U979 ( .A(KEYINPUT114), .B(n880), .ZN(n887) );
  NAND2_X1 U980 ( .A1(G115), .A2(n881), .ZN(n884) );
  NAND2_X1 U981 ( .A1(G127), .A2(n882), .ZN(n883) );
  NAND2_X1 U982 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U983 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U984 ( .A1(n887), .A2(n886), .ZN(n1002) );
  XOR2_X1 U985 ( .A(G160), .B(G162), .Z(n888) );
  XNOR2_X1 U986 ( .A(n993), .B(n888), .ZN(n889) );
  XNOR2_X1 U987 ( .A(n1002), .B(n889), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n890), .B(G164), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n897) );
  XNOR2_X1 U991 ( .A(n895), .B(KEYINPUT48), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n899) );
  XOR2_X1 U993 ( .A(n899), .B(n898), .Z(n900) );
  NOR2_X1 U994 ( .A1(G37), .A2(n900), .ZN(G395) );
  XOR2_X1 U995 ( .A(KEYINPUT115), .B(n901), .Z(n903) );
  XNOR2_X1 U996 ( .A(n971), .B(G286), .ZN(n902) );
  XNOR2_X1 U997 ( .A(n903), .B(n902), .ZN(n905) );
  XNOR2_X1 U998 ( .A(n964), .B(G301), .ZN(n904) );
  XNOR2_X1 U999 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n906), .ZN(G397) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n907) );
  XOR2_X1 U1002 ( .A(KEYINPUT49), .B(n907), .Z(n910) );
  NOR2_X1 U1003 ( .A1(G401), .A2(n914), .ZN(n908) );
  XNOR2_X1 U1004 ( .A(KEYINPUT116), .B(n908), .ZN(n909) );
  NAND2_X1 U1005 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1006 ( .A(KEYINPUT117), .B(n911), .ZN(n913) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(n913), .A2(n912), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(n914), .ZN(G319) );
  INV_X1 U1011 ( .A(G69), .ZN(G235) );
  INV_X1 U1012 ( .A(n915), .ZN(G223) );
  INV_X1 U1013 ( .A(G301), .ZN(G171) );
  INV_X1 U1014 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U1015 ( .A(G1966), .B(G21), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(G5), .B(G1961), .ZN(n916) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n927) );
  XOR2_X1 U1018 ( .A(G1348), .B(KEYINPUT59), .Z(n918) );
  XNOR2_X1 U1019 ( .A(G4), .B(n918), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(G20), .B(G1956), .ZN(n919) );
  NOR2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(G1341), .B(G19), .ZN(n922) );
  XNOR2_X1 U1023 ( .A(G1981), .B(G6), .ZN(n921) );
  NOR2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  XOR2_X1 U1026 ( .A(KEYINPUT60), .B(n925), .Z(n926) );
  NAND2_X1 U1027 ( .A1(n927), .A2(n926), .ZN(n934) );
  XNOR2_X1 U1028 ( .A(G1971), .B(G22), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(G23), .B(G1976), .ZN(n928) );
  NOR2_X1 U1030 ( .A1(n929), .A2(n928), .ZN(n931) );
  XOR2_X1 U1031 ( .A(G1986), .B(G24), .Z(n930) );
  NAND2_X1 U1032 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(KEYINPUT58), .B(n932), .ZN(n933) );
  NOR2_X1 U1034 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(n935), .B(KEYINPUT61), .ZN(n937) );
  XNOR2_X1 U1036 ( .A(G16), .B(KEYINPUT127), .ZN(n936) );
  NAND2_X1 U1037 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1038 ( .A1(G11), .A2(n938), .ZN(n1018) );
  INV_X1 U1039 ( .A(G29), .ZN(n1011) );
  XOR2_X1 U1040 ( .A(n1011), .B(KEYINPUT125), .Z(n962) );
  XNOR2_X1 U1041 ( .A(G2084), .B(G34), .ZN(n939) );
  XNOR2_X1 U1042 ( .A(n939), .B(KEYINPUT54), .ZN(n958) );
  XNOR2_X1 U1043 ( .A(KEYINPUT122), .B(KEYINPUT53), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(KEYINPUT121), .B(G2072), .ZN(n940) );
  XNOR2_X1 U1045 ( .A(n940), .B(G33), .ZN(n947) );
  XOR2_X1 U1046 ( .A(G2067), .B(G26), .Z(n942) );
  XOR2_X1 U1047 ( .A(G1996), .B(G32), .Z(n941) );
  NAND2_X1 U1048 ( .A1(n942), .A2(n941), .ZN(n945) );
  XNOR2_X1 U1049 ( .A(G27), .B(n943), .ZN(n944) );
  NOR2_X1 U1050 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1051 ( .A1(n947), .A2(n946), .ZN(n950) );
  XOR2_X1 U1052 ( .A(G1991), .B(G25), .Z(n948) );
  NAND2_X1 U1053 ( .A1(G28), .A2(n948), .ZN(n949) );
  NOR2_X1 U1054 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1055 ( .A(n952), .B(n951), .ZN(n955) );
  XNOR2_X1 U1056 ( .A(G2090), .B(G35), .ZN(n953) );
  XNOR2_X1 U1057 ( .A(KEYINPUT120), .B(n953), .ZN(n954) );
  NOR2_X1 U1058 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1059 ( .A(n956), .B(KEYINPUT123), .ZN(n957) );
  NOR2_X1 U1060 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1061 ( .A(n959), .B(KEYINPUT124), .ZN(n960) );
  XNOR2_X1 U1062 ( .A(n960), .B(KEYINPUT55), .ZN(n961) );
  NAND2_X1 U1063 ( .A1(n962), .A2(n961), .ZN(n1016) );
  XOR2_X1 U1064 ( .A(KEYINPUT56), .B(G16), .Z(n987) );
  XNOR2_X1 U1065 ( .A(n963), .B(KEYINPUT126), .ZN(n968) );
  XOR2_X1 U1066 ( .A(G171), .B(G1961), .Z(n966) );
  XNOR2_X1 U1067 ( .A(n964), .B(G1341), .ZN(n965) );
  NOR2_X1 U1068 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1069 ( .A1(n968), .A2(n967), .ZN(n985) );
  NAND2_X1 U1070 ( .A1(n970), .A2(n969), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(n971), .B(G1348), .ZN(n976) );
  XOR2_X1 U1072 ( .A(G166), .B(G1971), .Z(n974) );
  XNOR2_X1 U1073 ( .A(n972), .B(G1956), .ZN(n973) );
  NOR2_X1 U1074 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1075 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1076 ( .A1(n978), .A2(n977), .ZN(n983) );
  XOR2_X1 U1077 ( .A(G168), .B(G1966), .Z(n979) );
  NOR2_X1 U1078 ( .A1(n980), .A2(n979), .ZN(n981) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n981), .Z(n982) );
  NAND2_X1 U1080 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1081 ( .A1(n985), .A2(n984), .ZN(n986) );
  NOR2_X1 U1082 ( .A1(n987), .A2(n986), .ZN(n1014) );
  XOR2_X1 U1083 ( .A(G2090), .B(G162), .Z(n988) );
  NOR2_X1 U1084 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1085 ( .A(KEYINPUT51), .B(n990), .Z(n992) );
  NAND2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n999) );
  XNOR2_X1 U1087 ( .A(G160), .B(G2084), .ZN(n994) );
  NAND2_X1 U1088 ( .A1(n994), .A2(n993), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1090 ( .A(KEYINPUT118), .B(n997), .Z(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1007) );
  XOR2_X1 U1093 ( .A(G2072), .B(n1002), .Z(n1004) );
  XOR2_X1 U1094 ( .A(G164), .B(G2078), .Z(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1096 ( .A(KEYINPUT50), .B(n1005), .Z(n1006) );
  NOR2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XOR2_X1 U1098 ( .A(KEYINPUT52), .B(n1008), .Z(n1009) );
  NOR2_X1 U1099 ( .A1(KEYINPUT55), .A2(n1009), .ZN(n1010) );
  NOR2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1101 ( .A(KEYINPUT119), .B(n1012), .Z(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1105 ( .A(KEYINPUT62), .B(n1019), .Z(G150) );
  INV_X1 U1106 ( .A(G150), .ZN(G311) );
endmodule

