//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 1 0 0 1 0 0 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:41 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n577, new_n578, new_n579, new_n580, new_n581, new_n582,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n633, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT64), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(G234));
  NAND2_X1  g024(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  XNOR2_X1  g030(.A(G325), .B(KEYINPUT66), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI211_X1 g038(.A(G137), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n461), .A2(G101), .A3(G2104), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n465), .B1(new_n464), .B2(new_n466), .ZN(new_n468));
  OR2_X1    g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OR2_X1    g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AND2_X1   g048(.A1(G113), .A2(G2104), .ZN(new_n474));
  OAI21_X1  g049(.A(G2105), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n469), .A2(new_n475), .ZN(G160));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(G112), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n477), .B1(new_n478), .B2(G2105), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n462), .A2(new_n463), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n461), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n479), .B1(new_n481), .B2(G124), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT68), .B1(new_n480), .B2(G2105), .ZN(new_n483));
  XNOR2_X1  g058(.A(KEYINPUT3), .B(G2104), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT68), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n484), .A2(new_n485), .A3(new_n461), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(G136), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n482), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G162));
  NAND2_X1  g065(.A1(G126), .A2(G2105), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n471), .B2(new_n472), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n461), .A2(G114), .ZN(new_n493));
  OAI21_X1  g068(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT69), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n497), .A2(new_n499), .A3(G2104), .ZN(new_n500));
  AND2_X1   g075(.A1(G126), .A2(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n501), .B1(new_n462), .B2(new_n463), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n500), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  OAI211_X1 g079(.A(G138), .B(new_n461), .C1(new_n462), .C2(new_n463), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n484), .A2(new_n507), .A3(G138), .A4(new_n461), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n496), .A2(new_n504), .B1(new_n506), .B2(new_n508), .ZN(G164));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  OAI21_X1  g085(.A(KEYINPUT71), .B1(new_n510), .B2(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n512), .A2(new_n513), .A3(G543), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n511), .A2(new_n514), .B1(KEYINPUT5), .B2(new_n510), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  OAI211_X1 g096(.A(G50), .B(G543), .C1(new_n520), .C2(new_n521), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n522), .A2(KEYINPUT70), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(KEYINPUT70), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(KEYINPUT6), .A2(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n515), .A2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G88), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n519), .A2(new_n525), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(G166));
  NAND3_X1  g108(.A1(new_n515), .A2(G89), .A3(new_n528), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n510), .B1(new_n526), .B2(new_n527), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(KEYINPUT7), .ZN(new_n538));
  AOI22_X1  g113(.A1(G51), .A2(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AND2_X1   g114(.A1(G63), .A2(G651), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n515), .A2(KEYINPUT72), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(KEYINPUT72), .B1(new_n515), .B2(new_n540), .ZN(new_n542));
  OAI211_X1 g117(.A(new_n534), .B(new_n539), .C1(new_n541), .C2(new_n542), .ZN(G286));
  INV_X1    g118(.A(G286), .ZN(G168));
  NAND2_X1  g119(.A1(new_n535), .A2(G52), .ZN(new_n545));
  XOR2_X1   g120(.A(KEYINPUT73), .B(G90), .Z(new_n546));
  NAND3_X1  g121(.A1(new_n515), .A2(new_n528), .A3(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G651), .ZN(new_n549));
  OAI211_X1 g124(.A(new_n545), .B(new_n547), .C1(new_n548), .C2(new_n549), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  AOI22_X1  g126(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n552), .A2(new_n549), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n515), .A2(G81), .A3(new_n528), .ZN(new_n554));
  XOR2_X1   g129(.A(KEYINPUT74), .B(G43), .Z(new_n555));
  NAND2_X1  g130(.A1(new_n535), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT75), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n554), .A2(new_n559), .A3(new_n556), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n553), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT76), .ZN(G188));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  AND3_X1   g143(.A1(new_n535), .A2(new_n568), .A3(G53), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n568), .B1(new_n535), .B2(G53), .ZN(new_n570));
  INV_X1    g145(.A(G91), .ZN(new_n571));
  OAI22_X1  g146(.A1(new_n569), .A2(new_n570), .B1(new_n529), .B2(new_n571), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n515), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n573), .A2(new_n549), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G299));
  INV_X1    g151(.A(KEYINPUT77), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n519), .A2(new_n525), .A3(new_n531), .A4(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(G88), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n523), .A2(new_n524), .B1(new_n529), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n549), .B1(new_n516), .B2(new_n517), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT77), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g157(.A1(new_n578), .A2(new_n582), .ZN(G303));
  OAI21_X1  g158(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n515), .A2(G87), .A3(new_n528), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n535), .A2(G49), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT78), .A4(new_n586), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G288));
  OAI211_X1 g167(.A(G48), .B(G543), .C1(new_n520), .C2(new_n521), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT79), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n535), .A2(new_n595), .A3(G48), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n530), .A2(G86), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n515), .A2(G61), .ZN(new_n598));
  NAND2_X1  g173(.A1(G73), .A2(G543), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n549), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT80), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n597), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G86), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n595), .B1(new_n535), .B2(G48), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n593), .A2(KEYINPUT79), .ZN(new_n606));
  OAI22_X1  g181(.A1(new_n604), .A2(new_n529), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(KEYINPUT80), .B1(new_n607), .B2(new_n600), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n603), .A2(new_n608), .ZN(G305));
  AND2_X1   g184(.A1(G72), .A2(G543), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n515), .B2(G60), .ZN(new_n611));
  OR3_X1    g186(.A1(new_n611), .A2(KEYINPUT81), .A3(new_n549), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n530), .A2(G85), .B1(G47), .B2(new_n535), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT81), .B1(new_n611), .B2(new_n549), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(G290));
  NAND2_X1  g190(.A1(G301), .A2(G868), .ZN(new_n616));
  INV_X1    g191(.A(G92), .ZN(new_n617));
  OAI21_X1  g192(.A(KEYINPUT82), .B1(new_n529), .B2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n619));
  NAND4_X1  g194(.A1(new_n515), .A2(new_n619), .A3(G92), .A4(new_n528), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT10), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n535), .A2(G54), .ZN(new_n624));
  AOI22_X1  g199(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(new_n549), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n618), .A2(KEYINPUT10), .A3(new_n620), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n623), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n616), .B1(new_n630), .B2(G868), .ZN(G284));
  OAI21_X1  g206(.A(new_n616), .B1(new_n630), .B2(G868), .ZN(G321));
  NAND2_X1  g207(.A1(G286), .A2(G868), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n633), .B1(new_n575), .B2(G868), .ZN(G297));
  OAI21_X1  g209(.A(new_n633), .B1(new_n575), .B2(G868), .ZN(G280));
  INV_X1    g210(.A(G559), .ZN(new_n636));
  OAI21_X1  g211(.A(new_n630), .B1(new_n636), .B2(G860), .ZN(G148));
  INV_X1    g212(.A(new_n561), .ZN(new_n638));
  INV_X1    g213(.A(G868), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n629), .A2(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n641), .B2(new_n639), .ZN(G323));
  XNOR2_X1  g217(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OAI21_X1  g218(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n644));
  INV_X1    g219(.A(G111), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n644), .B1(new_n645), .B2(G2105), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n481), .B2(G123), .ZN(new_n647));
  INV_X1    g222(.A(G135), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n647), .B1(new_n487), .B2(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(new_n649), .B(KEYINPUT83), .Z(new_n650));
  OR2_X1    g225(.A1(new_n650), .A2(G2096), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(G2096), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n461), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n653), .B(KEYINPUT12), .Z(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT13), .ZN(new_n655));
  XOR2_X1   g230(.A(new_n655), .B(G2100), .Z(new_n656));
  NAND3_X1  g231(.A1(new_n651), .A2(new_n652), .A3(new_n656), .ZN(G156));
  XOR2_X1   g232(.A(G2443), .B(G2446), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT85), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(G2451), .ZN(new_n660));
  XOR2_X1   g235(.A(G1341), .B(G1348), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2427), .B(G2438), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2430), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT15), .B(G2435), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n664), .A2(new_n665), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n667), .A3(KEYINPUT14), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n662), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G2454), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G14), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n669), .A2(new_n671), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(G401));
  XOR2_X1   g250(.A(G2072), .B(G2078), .Z(new_n676));
  AND2_X1   g251(.A1(new_n676), .A2(KEYINPUT87), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  XNOR2_X1  g253(.A(G2067), .B(G2678), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(KEYINPUT87), .B2(new_n676), .ZN(new_n681));
  OR2_X1    g256(.A1(new_n676), .A2(KEYINPUT17), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n676), .A2(KEYINPUT17), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n682), .B(new_n683), .C1(new_n678), .C2(new_n679), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n678), .A2(new_n679), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n676), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT86), .B(KEYINPUT18), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(G2096), .B(G2100), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(G227));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  INV_X1    g268(.A(KEYINPUT19), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(G1956), .B(G2474), .Z(new_n696));
  XOR2_X1   g271(.A(G1961), .B(G1966), .Z(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n700));
  XOR2_X1   g275(.A(new_n699), .B(new_n700), .Z(new_n701));
  NOR2_X1   g276(.A1(new_n696), .A2(new_n697), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n695), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT89), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n695), .A2(new_n698), .A3(new_n702), .ZN(new_n705));
  NOR3_X1   g280(.A1(new_n701), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XOR2_X1   g283(.A(G1991), .B(G1996), .Z(new_n709));
  XOR2_X1   g284(.A(new_n708), .B(new_n709), .Z(new_n710));
  XNOR2_X1  g285(.A(G1981), .B(G1986), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n708), .B(new_n709), .ZN(new_n713));
  INV_X1    g288(.A(new_n711), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n712), .A2(new_n715), .ZN(G229));
  XNOR2_X1  g291(.A(KEYINPUT90), .B(G16), .ZN(new_n717));
  MUX2_X1   g292(.A(new_n532), .B(G22), .S(new_n717), .Z(new_n718));
  INV_X1    g293(.A(G1971), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(G305), .A2(G16), .ZN(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n722), .A2(G6), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(KEYINPUT32), .B(G1981), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g301(.A(new_n725), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n721), .A2(new_n727), .A3(new_n723), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n722), .A2(G23), .ZN(new_n729));
  INV_X1    g304(.A(new_n587), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(new_n722), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT33), .B(G1976), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND4_X1  g308(.A1(new_n720), .A2(new_n726), .A3(new_n728), .A4(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n734), .A2(KEYINPUT34), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  MUX2_X1   g311(.A(G290), .B(G24), .S(new_n717), .Z(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(G1986), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G25), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n483), .A2(new_n486), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G131), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n743));
  INV_X1    g318(.A(G107), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n743), .B1(new_n744), .B2(G2105), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n481), .B2(G119), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n742), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n740), .B1(new_n748), .B2(new_n739), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT35), .B(G1991), .Z(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n749), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n738), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(new_n734), .B2(KEYINPUT34), .ZN(new_n754));
  OAI21_X1  g329(.A(KEYINPUT36), .B1(new_n736), .B2(new_n754), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n734), .A2(KEYINPUT34), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT36), .ZN(new_n757));
  NAND4_X1  g332(.A1(new_n756), .A2(new_n735), .A3(new_n757), .A4(new_n753), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n650), .A2(new_n739), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT31), .B(G11), .ZN(new_n761));
  XNOR2_X1  g336(.A(KEYINPUT97), .B(G28), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(KEYINPUT30), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n762), .A2(KEYINPUT30), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(new_n739), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT91), .B(KEYINPUT28), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n739), .A2(G26), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n483), .A2(G140), .A3(new_n486), .ZN(new_n770));
  OAI21_X1  g345(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n771));
  INV_X1    g346(.A(G116), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n771), .B1(new_n772), .B2(G2105), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n481), .B2(G128), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n769), .B1(new_n776), .B2(new_n739), .ZN(new_n777));
  OAI221_X1 g352(.A(new_n761), .B1(new_n763), .B2(new_n765), .C1(new_n777), .C2(G2067), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n777), .A2(G2067), .ZN(new_n779));
  NOR3_X1   g354(.A1(new_n760), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n739), .A2(G27), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G164), .B2(new_n739), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G2078), .ZN(new_n783));
  AND2_X1   g358(.A1(new_n739), .A2(G32), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n741), .A2(G141), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n481), .A2(G129), .ZN(new_n786));
  NAND3_X1  g361(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT26), .Z(new_n788));
  NAND3_X1  g363(.A1(new_n461), .A2(G105), .A3(G2104), .ZN(new_n789));
  AND3_X1   g364(.A1(new_n786), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n785), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n784), .B1(new_n791), .B2(G29), .ZN(new_n792));
  XOR2_X1   g367(.A(KEYINPUT27), .B(G1996), .Z(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT96), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n792), .A2(new_n795), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n783), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n739), .A2(G35), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(G162), .B2(new_n739), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n800), .A2(KEYINPUT29), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n800), .A2(KEYINPUT29), .ZN(new_n802));
  OR3_X1    g377(.A1(new_n801), .A2(new_n802), .A3(G2090), .ZN(new_n803));
  INV_X1    g378(.A(G34), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n804), .A2(KEYINPUT24), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(KEYINPUT24), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n739), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G160), .B2(new_n739), .ZN(new_n808));
  INV_X1    g383(.A(G2084), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n808), .B(new_n809), .ZN(new_n810));
  NAND4_X1  g385(.A1(new_n780), .A2(new_n798), .A3(new_n803), .A4(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n717), .A2(G20), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT23), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(new_n575), .B2(new_n722), .ZN(new_n814));
  INV_X1    g389(.A(G1956), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(G2090), .B1(new_n801), .B2(new_n802), .ZN(new_n817));
  AOI21_X1  g392(.A(KEYINPUT99), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n811), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(G115), .A2(G2104), .ZN(new_n820));
  INV_X1    g395(.A(G127), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n820), .B1(new_n480), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT92), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT92), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(new_n820), .C1(new_n480), .C2(new_n821), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n823), .A2(new_n825), .A3(G2105), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n483), .A2(G139), .A3(new_n486), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT25), .Z(new_n829));
  NAND3_X1  g404(.A1(new_n826), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n830), .A2(KEYINPUT93), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(KEYINPUT93), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n739), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n739), .A2(G33), .ZN(new_n834));
  OR3_X1    g409(.A1(new_n833), .A2(KEYINPUT94), .A3(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(G2072), .ZN(new_n836));
  OAI21_X1  g411(.A(KEYINPUT94), .B1(new_n833), .B2(new_n834), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n717), .A2(G19), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n561), .B2(new_n717), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(G1341), .ZN(new_n841));
  AND2_X1   g416(.A1(new_n722), .A2(G5), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(G301), .B2(G16), .ZN(new_n843));
  INV_X1    g418(.A(G1961), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT98), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n722), .A2(G21), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(G168), .B2(new_n722), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n848), .A2(G1966), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(G1966), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n843), .A2(new_n844), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR4_X1   g427(.A1(new_n841), .A2(new_n846), .A3(new_n849), .A4(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n819), .A2(new_n838), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT95), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n835), .A2(new_n837), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n855), .B1(new_n856), .B2(G2072), .ZN(new_n857));
  AOI211_X1 g432(.A(KEYINPUT95), .B(new_n836), .C1(new_n835), .C2(new_n837), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n630), .A2(G16), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n860), .B1(G4), .B2(G16), .ZN(new_n861));
  INV_X1    g436(.A(G1348), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n816), .A2(new_n817), .A3(KEYINPUT99), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NOR3_X1   g441(.A1(new_n854), .A2(new_n859), .A3(new_n866), .ZN(new_n867));
  AND3_X1   g442(.A1(new_n759), .A2(new_n867), .A3(KEYINPUT100), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT100), .B1(new_n759), .B2(new_n867), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(new_n869), .ZN(G311));
  NAND2_X1  g445(.A1(new_n759), .A2(new_n867), .ZN(G150));
  NAND2_X1  g446(.A1(new_n630), .A2(G559), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT38), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n874));
  AND2_X1   g449(.A1(G80), .A2(G543), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n875), .B1(new_n515), .B2(G67), .ZN(new_n876));
  OAI21_X1  g451(.A(G651), .B1(new_n876), .B2(KEYINPUT101), .ZN(new_n877));
  INV_X1    g452(.A(G67), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n513), .A2(G543), .ZN(new_n879));
  AOI211_X1 g454(.A(new_n878), .B(new_n879), .C1(new_n511), .C2(new_n514), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n881));
  NOR3_X1   g456(.A1(new_n880), .A2(new_n881), .A3(new_n875), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n874), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n876), .A2(KEYINPUT101), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n881), .B1(new_n880), .B2(new_n875), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT102), .A4(G651), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n535), .A2(G55), .ZN(new_n887));
  INV_X1    g462(.A(G93), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n887), .B1(new_n529), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n883), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n891), .A2(new_n638), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n884), .A2(new_n885), .A3(G651), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n889), .B1(new_n893), .B2(new_n874), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n894), .A2(new_n561), .A3(new_n886), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n873), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT39), .ZN(new_n898));
  AOI21_X1  g473(.A(G860), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n899), .B1(new_n898), .B2(new_n897), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n891), .A2(G860), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(KEYINPUT37), .Z(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(G145));
  NAND3_X1  g478(.A1(new_n741), .A2(KEYINPUT103), .A3(G142), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  INV_X1    g480(.A(G142), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n905), .B1(new_n487), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT104), .ZN(new_n910));
  INV_X1    g485(.A(G118), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n909), .A2(new_n910), .B1(new_n911), .B2(G2105), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(new_n910), .B2(new_n909), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n481), .A2(G130), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n908), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n742), .A2(KEYINPUT105), .A3(new_n746), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(KEYINPUT105), .B1(new_n742), .B2(new_n746), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n918), .A2(new_n919), .A3(new_n654), .ZN(new_n920));
  INV_X1    g495(.A(new_n654), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT105), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n747), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n921), .B1(new_n923), .B2(new_n917), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n916), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n654), .B1(new_n918), .B2(new_n919), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n923), .A2(new_n921), .A3(new_n917), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n926), .A2(new_n927), .A3(new_n915), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n831), .A2(new_n832), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n791), .A2(new_n775), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n776), .A2(new_n785), .A3(new_n790), .ZN(new_n933));
  AND2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n500), .A2(new_n502), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n936), .B1(new_n506), .B2(new_n508), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n932), .A2(new_n933), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n938), .A2(new_n832), .A3(new_n831), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n935), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n937), .B1(new_n935), .B2(new_n939), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n930), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n935), .A2(new_n939), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n506), .A2(new_n508), .ZN(new_n945));
  INV_X1    g520(.A(new_n936), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n944), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n948), .A2(new_n929), .A3(new_n940), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n943), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(G160), .B(new_n489), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(new_n650), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT106), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n950), .A2(KEYINPUT106), .A3(new_n953), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n943), .B(new_n952), .C1(new_n949), .C2(KEYINPUT107), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n949), .A2(KEYINPUT107), .ZN(new_n961));
  AOI21_X1  g536(.A(G37), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n958), .A2(new_n962), .A3(KEYINPUT40), .ZN(new_n963));
  AOI21_X1  g538(.A(KEYINPUT40), .B1(new_n958), .B2(new_n962), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n963), .A2(new_n964), .ZN(G395));
  NAND2_X1  g540(.A1(new_n891), .A2(new_n639), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT41), .ZN(new_n967));
  AND4_X1   g542(.A1(new_n575), .A2(new_n623), .A3(new_n628), .A4(new_n627), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n626), .B1(new_n621), .B2(new_n622), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n575), .B1(new_n969), .B2(new_n628), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n967), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n629), .A2(G299), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n575), .A3(new_n628), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n972), .A2(KEYINPUT41), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n892), .B2(new_n895), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n892), .A2(new_n895), .A3(new_n976), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n641), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n979), .ZN(new_n981));
  INV_X1    g556(.A(new_n641), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n981), .A2(new_n977), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n975), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n978), .A2(new_n641), .A3(new_n979), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n982), .B1(new_n981), .B2(new_n977), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT109), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n987), .B1(new_n968), .B2(new_n970), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n972), .A2(KEYINPUT109), .A3(new_n973), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n985), .A2(new_n986), .A3(new_n988), .A4(new_n989), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n984), .A2(KEYINPUT111), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT111), .B1(new_n984), .B2(new_n990), .ZN(new_n992));
  NAND2_X1  g567(.A1(G290), .A2(new_n730), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n612), .A2(new_n587), .A3(new_n613), .A4(new_n614), .ZN(new_n994));
  AND3_X1   g569(.A1(new_n993), .A2(G166), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(G166), .B1(new_n993), .B2(new_n994), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n997), .B1(new_n603), .B2(new_n608), .ZN(new_n998));
  AND3_X1   g573(.A1(new_n603), .A2(new_n608), .A3(new_n997), .ZN(new_n999));
  OAI22_X1  g574(.A1(new_n995), .A2(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n993), .A2(new_n994), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(new_n532), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n999), .A2(new_n998), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n993), .A2(G166), .A3(new_n994), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT42), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n991), .B1(new_n992), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1007), .ZN(new_n1009));
  NAND4_X1  g584(.A1(new_n1009), .A2(KEYINPUT111), .A3(new_n984), .A4(new_n990), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n966), .B1(new_n1011), .B2(new_n639), .ZN(G295));
  OAI21_X1  g587(.A(new_n966), .B1(new_n1011), .B2(new_n639), .ZN(G331));
  INV_X1    g588(.A(KEYINPUT44), .ZN(new_n1014));
  AND2_X1   g589(.A1(new_n1000), .A2(new_n1005), .ZN(new_n1015));
  XNOR2_X1  g590(.A(G286), .B(G301), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n561), .B1(new_n894), .B2(new_n886), .ZN(new_n1018));
  AND4_X1   g593(.A1(new_n561), .A2(new_n883), .A3(new_n886), .A4(new_n890), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n892), .A2(new_n895), .A3(new_n1016), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1020), .A2(new_n971), .A3(new_n974), .A4(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1020), .A2(new_n1021), .B1(new_n988), .B2(new_n989), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1015), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT43), .ZN(new_n1026));
  INV_X1    g601(.A(G37), .ZN(new_n1027));
  NOR2_X1   g602(.A1(new_n968), .A2(new_n970), .ZN(new_n1028));
  AND3_X1   g603(.A1(new_n892), .A2(new_n895), .A3(new_n1016), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1016), .B1(new_n892), .B2(new_n895), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1006), .A2(new_n1031), .A3(new_n1022), .ZN(new_n1032));
  NAND4_X1  g607(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .A4(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(KEYINPUT113), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1032), .A2(new_n1027), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT113), .ZN(new_n1036));
  NAND4_X1  g611(.A1(new_n1035), .A2(new_n1036), .A3(new_n1026), .A4(new_n1025), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1032), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1031), .A2(new_n1022), .ZN(new_n1040));
  AOI21_X1  g615(.A(G37), .B1(new_n1040), .B2(new_n1015), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1039), .B1(new_n1041), .B2(KEYINPUT112), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT112), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1006), .B1(new_n1022), .B2(new_n1031), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(new_n1044), .B2(G37), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1026), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1014), .B1(new_n1038), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(KEYINPUT43), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1048));
  AND3_X1   g623(.A1(new_n1035), .A2(KEYINPUT43), .A3(new_n1025), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT44), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1047), .A2(new_n1050), .ZN(G397));
  INV_X1    g626(.A(G1384), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n947), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT114), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT45), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI211_X1 g630(.A(G40), .B(new_n475), .C1(new_n467), .C2(new_n468), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n937), .A2(G1384), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(KEYINPUT114), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1055), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n748), .A2(new_n750), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n747), .A2(new_n751), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  XNOR2_X1  g639(.A(new_n775), .B(G2067), .ZN(new_n1065));
  AND2_X1   g640(.A1(new_n791), .A2(G1996), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1061), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  OR2_X1    g642(.A1(new_n1060), .A2(G1996), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(new_n791), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT115), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1068), .A2(KEYINPUT115), .A3(new_n791), .ZN(new_n1072));
  OAI211_X1 g647(.A(new_n1064), .B(new_n1067), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1073));
  XNOR2_X1  g648(.A(G290), .B(G1986), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1073), .B1(new_n1061), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT123), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT116), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n1077), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT50), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n947), .A2(new_n1079), .A3(new_n1052), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(new_n1057), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(new_n504), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n503), .B1(new_n500), .B2(new_n502), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n945), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(new_n1052), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1077), .B1(new_n1085), .B2(KEYINPUT50), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1076), .B1(new_n1081), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(G164), .A2(G1384), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT116), .B1(new_n1088), .B2(new_n1079), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1056), .B1(new_n1058), .B2(new_n1079), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1089), .A2(KEYINPUT123), .A3(new_n1078), .A4(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1087), .A2(new_n844), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT45), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n937), .B2(G1384), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1093), .B1(new_n1057), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1088), .A2(KEYINPUT45), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1057), .A2(new_n1095), .A3(new_n1093), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1100), .A2(G2078), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1097), .A2(new_n1098), .A3(new_n1099), .A4(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1085), .A2(new_n1094), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1056), .B1(new_n1058), .B2(KEYINPUT45), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1100), .B1(new_n1105), .B2(G2078), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1092), .A2(new_n1102), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(G171), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1055), .A2(new_n1059), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1109), .A2(new_n1104), .A3(new_n1101), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1092), .A2(G301), .A3(new_n1106), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1108), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1105), .A2(new_n719), .ZN(new_n1115));
  INV_X1    g690(.A(G2090), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1089), .A2(new_n1116), .A3(new_n1078), .A4(new_n1090), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1117), .A3(KEYINPUT117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(G8), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n578), .A2(new_n582), .A3(G8), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n1121));
  XNOR2_X1  g696(.A(new_n1120), .B(new_n1121), .ZN(new_n1122));
  AOI21_X1  g697(.A(KEYINPUT117), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1119), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT49), .ZN(new_n1125));
  INV_X1    g700(.A(G1981), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1126), .B1(new_n597), .B2(new_n601), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n607), .A2(new_n600), .A3(G1981), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g704(.A(G8), .B1(new_n1053), .B2(new_n1056), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n597), .A2(new_n601), .A3(new_n1126), .ZN(new_n1132));
  OAI21_X1  g707(.A(G1981), .B1(new_n607), .B2(new_n600), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1132), .A2(new_n1133), .A3(KEYINPUT49), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1129), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n584), .A2(new_n585), .A3(G1976), .A4(new_n586), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1136), .B(KEYINPUT119), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT52), .ZN(new_n1138));
  INV_X1    g713(.A(G1976), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n589), .A2(new_n1139), .A3(new_n590), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1131), .A2(new_n1137), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n1142));
  XNOR2_X1  g717(.A(new_n1136), .B(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(KEYINPUT52), .B1(new_n1143), .B2(new_n1130), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1135), .A2(new_n1141), .A3(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1084), .A2(new_n1079), .A3(new_n1052), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT50), .B1(new_n937), .B2(G1384), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1146), .A2(new_n1057), .A3(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(G2090), .ZN(new_n1149));
  AOI21_X1  g724(.A(G1971), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1150));
  OAI21_X1  g725(.A(G8), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1122), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1145), .A2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n1124), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(G1966), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1099), .A2(new_n1098), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1155), .B1(new_n1156), .B2(new_n1096), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1089), .A2(new_n809), .A3(new_n1078), .A4(new_n1090), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1157), .A2(G168), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(G8), .ZN(new_n1160));
  AOI21_X1  g735(.A(G168), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT51), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT51), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1159), .A2(new_n1163), .A3(G8), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND4_X1  g740(.A1(new_n1092), .A2(new_n1102), .A3(G301), .A4(new_n1106), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1092), .A2(new_n1106), .A3(new_n1110), .ZN(new_n1167));
  OAI211_X1 g742(.A(KEYINPUT54), .B(new_n1166), .C1(new_n1167), .C2(G301), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1114), .A2(new_n1154), .A3(new_n1165), .A4(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(KEYINPUT58), .B(G1341), .ZN(new_n1172));
  OAI22_X1  g747(.A1(new_n1105), .A2(G1996), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(KEYINPUT125), .A2(KEYINPUT59), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n561), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1173), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g752(.A1(KEYINPUT125), .A2(KEYINPUT59), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n1177), .B(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n575), .B(KEYINPUT57), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1148), .A2(new_n815), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(KEYINPUT121), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT121), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1148), .A2(new_n1183), .A3(new_n815), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1182), .A2(new_n1184), .ZN(new_n1185));
  XNOR2_X1  g760(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(G2072), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1103), .A2(new_n1104), .A3(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1180), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n1190));
  AOI21_X1  g765(.A(KEYINPUT61), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1184), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1183), .B1(new_n1148), .B2(new_n815), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1188), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1180), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1194), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1185), .A2(new_n1180), .A3(new_n1188), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1196), .A2(new_n1197), .A3(KEYINPUT126), .ZN(new_n1198));
  AOI21_X1  g773(.A(new_n1179), .B1(new_n1191), .B2(new_n1198), .ZN(new_n1199));
  INV_X1    g774(.A(G2067), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1171), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1201), .B1(new_n1202), .B2(G1348), .ZN(new_n1203));
  INV_X1    g778(.A(new_n1203), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1204), .A2(KEYINPUT60), .A3(new_n629), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT124), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1196), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1189), .A2(KEYINPUT124), .ZN(new_n1208));
  NAND4_X1  g783(.A1(new_n1207), .A2(new_n1208), .A3(KEYINPUT61), .A4(new_n1197), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT60), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n629), .B1(new_n1203), .B2(new_n1210), .ZN(new_n1211));
  OAI21_X1  g786(.A(new_n1211), .B1(new_n1210), .B2(new_n1203), .ZN(new_n1212));
  NAND4_X1  g787(.A1(new_n1199), .A2(new_n1205), .A3(new_n1209), .A4(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1204), .A2(new_n629), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1197), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g791(.A(new_n1169), .B1(new_n1213), .B2(new_n1216), .ZN(new_n1217));
  INV_X1    g792(.A(KEYINPUT63), .ZN(new_n1218));
  INV_X1    g793(.A(G8), .ZN(new_n1219));
  AOI21_X1  g794(.A(new_n1219), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1220));
  INV_X1    g795(.A(new_n1220), .ZN(new_n1221));
  NAND4_X1  g796(.A1(new_n1135), .A2(G168), .A3(new_n1141), .A4(new_n1144), .ZN(new_n1222));
  NOR2_X1   g797(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  OAI21_X1  g798(.A(new_n1122), .B1(new_n1119), .B2(new_n1123), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1218), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  INV_X1    g800(.A(new_n1145), .ZN(new_n1226));
  NOR2_X1   g801(.A1(G286), .A2(KEYINPUT63), .ZN(new_n1227));
  NAND3_X1  g802(.A1(new_n1152), .A2(new_n1220), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1229));
  INV_X1    g804(.A(KEYINPUT117), .ZN(new_n1230));
  NAND2_X1  g805(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g806(.A(new_n1121), .ZN(new_n1232));
  XNOR2_X1  g807(.A(new_n1120), .B(new_n1232), .ZN(new_n1233));
  NAND4_X1  g808(.A1(new_n1231), .A2(G8), .A3(new_n1233), .A4(new_n1118), .ZN(new_n1234));
  AOI21_X1  g809(.A(new_n1226), .B1(new_n1228), .B2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1129), .A2(new_n1134), .ZN(new_n1236));
  NAND3_X1  g811(.A1(new_n1236), .A2(new_n1139), .A3(new_n591), .ZN(new_n1237));
  AOI21_X1  g812(.A(new_n1130), .B1(new_n1237), .B2(new_n1132), .ZN(new_n1238));
  NOR3_X1   g813(.A1(new_n1225), .A2(new_n1235), .A3(new_n1238), .ZN(new_n1239));
  NOR3_X1   g814(.A1(new_n1124), .A2(new_n1108), .A3(new_n1153), .ZN(new_n1240));
  INV_X1    g815(.A(new_n1164), .ZN(new_n1241));
  INV_X1    g816(.A(new_n1161), .ZN(new_n1242));
  NAND3_X1  g817(.A1(new_n1242), .A2(G8), .A3(new_n1159), .ZN(new_n1243));
  AOI21_X1  g818(.A(new_n1241), .B1(new_n1243), .B2(KEYINPUT51), .ZN(new_n1244));
  INV_X1    g819(.A(KEYINPUT62), .ZN(new_n1245));
  OAI21_X1  g820(.A(new_n1240), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NOR2_X1   g821(.A1(new_n1165), .A2(KEYINPUT62), .ZN(new_n1247));
  OAI21_X1  g822(.A(new_n1239), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g823(.A(new_n1075), .B1(new_n1217), .B2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g824(.A(new_n1063), .B(new_n1067), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1250));
  NOR2_X1   g825(.A1(new_n775), .A2(G2067), .ZN(new_n1251));
  INV_X1    g826(.A(new_n1251), .ZN(new_n1252));
  AOI21_X1  g827(.A(new_n1060), .B1(new_n1250), .B2(new_n1252), .ZN(new_n1253));
  INV_X1    g828(.A(new_n1253), .ZN(new_n1254));
  INV_X1    g829(.A(KEYINPUT127), .ZN(new_n1255));
  XNOR2_X1  g830(.A(new_n1068), .B(KEYINPUT46), .ZN(new_n1256));
  INV_X1    g831(.A(KEYINPUT47), .ZN(new_n1257));
  OAI21_X1  g832(.A(new_n1061), .B1(new_n791), .B2(new_n1065), .ZN(new_n1258));
  AND3_X1   g833(.A1(new_n1256), .A2(new_n1257), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g834(.A(new_n1257), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1260));
  OR2_X1    g835(.A1(new_n1259), .A2(new_n1260), .ZN(new_n1261));
  NOR3_X1   g836(.A1(new_n1060), .A2(G1986), .A3(G290), .ZN(new_n1262));
  XNOR2_X1  g837(.A(new_n1262), .B(KEYINPUT48), .ZN(new_n1263));
  OR2_X1    g838(.A1(new_n1073), .A2(new_n1263), .ZN(new_n1264));
  NAND4_X1  g839(.A1(new_n1254), .A2(new_n1255), .A3(new_n1261), .A4(new_n1264), .ZN(new_n1265));
  OAI22_X1  g840(.A1(new_n1259), .A2(new_n1260), .B1(new_n1073), .B2(new_n1263), .ZN(new_n1266));
  OAI21_X1  g841(.A(KEYINPUT127), .B1(new_n1266), .B2(new_n1253), .ZN(new_n1267));
  NAND2_X1  g842(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g843(.A1(new_n1249), .A2(new_n1268), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g844(.A1(new_n1038), .A2(new_n1046), .ZN(new_n1271));
  NOR2_X1   g845(.A1(G227), .A2(new_n459), .ZN(new_n1272));
  OAI21_X1  g846(.A(new_n1272), .B1(new_n673), .B2(new_n674), .ZN(new_n1273));
  AOI21_X1  g847(.A(new_n1273), .B1(new_n712), .B2(new_n715), .ZN(new_n1274));
  AOI21_X1  g848(.A(new_n952), .B1(new_n943), .B2(new_n949), .ZN(new_n1275));
  XNOR2_X1  g849(.A(new_n1275), .B(new_n955), .ZN(new_n1276));
  INV_X1    g850(.A(new_n961), .ZN(new_n1277));
  OAI21_X1  g851(.A(new_n1027), .B1(new_n959), .B2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g852(.A(new_n1274), .B1(new_n1276), .B2(new_n1278), .ZN(new_n1279));
  NOR2_X1   g853(.A1(new_n1271), .A2(new_n1279), .ZN(G308));
  OAI221_X1 g854(.A(new_n1274), .B1(new_n1276), .B2(new_n1278), .C1(new_n1038), .C2(new_n1046), .ZN(G225));
endmodule


