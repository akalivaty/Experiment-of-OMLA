//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:12 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n614, new_n616, new_n617, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT66), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  INV_X1    g033(.A(G125), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G113), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT67), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G113), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n463), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2105), .ZN(new_n471));
  AND2_X1   g046(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n472));
  OAI211_X1 g047(.A(G137), .B(new_n471), .C1(new_n472), .C2(new_n460), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n465), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G101), .ZN(new_n476));
  AND3_X1   g051(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n474), .B1(new_n473), .B2(new_n476), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n470), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  NOR2_X1   g055(.A1(new_n472), .A2(new_n460), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n471), .B1(new_n461), .B2(new_n462), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  OR2_X1    g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n471), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n483), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  OAI211_X1 g064(.A(G126), .B(G2105), .C1(new_n472), .C2(new_n460), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n496), .B1(new_n472), .B2(new_n460), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n496), .B(new_n499), .C1(new_n460), .C2(new_n472), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n494), .B1(new_n498), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT6), .A2(G651), .ZN(new_n504));
  OAI211_X1 g079(.A(G50), .B(G543), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  OAI22_X1  g082(.A1(new_n506), .A2(new_n507), .B1(new_n503), .B2(new_n504), .ZN(new_n508));
  INV_X1    g083(.A(G88), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n505), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  OAI21_X1  g086(.A(G62), .B1(new_n507), .B2(new_n506), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  AOI21_X1  g088(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n502), .B1(new_n510), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G62), .ZN(new_n516));
  OR2_X1    g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  AOI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n513), .ZN(new_n520));
  OAI21_X1  g095(.A(G651), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n503), .A2(new_n504), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n517), .A2(new_n518), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n522), .A2(G88), .A3(new_n523), .ZN(new_n524));
  NAND4_X1  g099(.A1(new_n521), .A2(new_n524), .A3(KEYINPUT69), .A4(new_n505), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n515), .A2(new_n525), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n522), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G51), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n523), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n522), .A2(G89), .ZN(new_n533));
  NAND2_X1  g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n531), .A2(new_n535), .ZN(G168));
  XNOR2_X1  g111(.A(KEYINPUT70), .B(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n529), .A2(new_n537), .B1(new_n538), .B2(new_n508), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n511), .ZN(new_n541));
  OR2_X1    g116(.A1(new_n539), .A2(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  INV_X1    g118(.A(G43), .ZN(new_n544));
  INV_X1    g119(.A(G81), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n529), .A2(new_n544), .B1(new_n545), .B2(new_n508), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n547), .A2(new_n511), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  NAND4_X1  g125(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  AND2_X1   g129(.A1(new_n522), .A2(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G53), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT9), .ZN(new_n557));
  INV_X1    g132(.A(G78), .ZN(new_n558));
  INV_X1    g133(.A(G543), .ZN(new_n559));
  OR3_X1    g134(.A1(new_n558), .A2(new_n559), .A3(KEYINPUT71), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT71), .B1(new_n558), .B2(new_n559), .ZN(new_n561));
  XNOR2_X1  g136(.A(KEYINPUT72), .B(G65), .ZN(new_n562));
  OAI211_X1 g137(.A(new_n560), .B(new_n561), .C1(new_n532), .C2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(new_n508), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n563), .A2(G651), .B1(G91), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n557), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G168), .ZN(G286));
  INV_X1    g142(.A(G166), .ZN(G303));
  NAND2_X1  g143(.A1(new_n555), .A2(G49), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n564), .A2(G87), .ZN(new_n570));
  OAI21_X1  g145(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  OAI211_X1 g147(.A(G48), .B(G543), .C1(new_n503), .C2(new_n504), .ZN(new_n573));
  INV_X1    g148(.A(G86), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n508), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT73), .ZN(new_n578));
  INV_X1    g153(.A(G61), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n517), .B2(new_n518), .ZN(new_n580));
  OAI21_X1  g155(.A(G651), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n576), .A2(new_n581), .ZN(G305));
  INV_X1    g157(.A(G47), .ZN(new_n583));
  XOR2_X1   g158(.A(KEYINPUT74), .B(G85), .Z(new_n584));
  OAI22_X1  g159(.A1(new_n529), .A2(new_n583), .B1(new_n508), .B2(new_n584), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n511), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n588), .ZN(G290));
  NAND2_X1  g164(.A1(G301), .A2(G868), .ZN(new_n590));
  OR2_X1    g165(.A1(new_n529), .A2(KEYINPUT76), .ZN(new_n591));
  INV_X1    g166(.A(G54), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n592), .B1(new_n529), .B2(KEYINPUT76), .ZN(new_n593));
  XOR2_X1   g168(.A(KEYINPUT75), .B(KEYINPUT10), .Z(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  OR3_X1    g170(.A1(new_n508), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n594), .B1(new_n508), .B2(new_n595), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n591), .A2(new_n593), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(KEYINPUT77), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(KEYINPUT77), .ZN(new_n601));
  AOI22_X1  g176(.A1(G66), .A2(new_n523), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT78), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n511), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(new_n603), .B2(new_n602), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n590), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n590), .B1(new_n607), .B2(G868), .ZN(G321));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(G299), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(new_n610), .B2(G168), .ZN(G297));
  OAI21_X1  g187(.A(new_n611), .B1(new_n610), .B2(G168), .ZN(G280));
  INV_X1    g188(.A(G559), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n607), .B1(new_n614), .B2(G860), .ZN(G148));
  NAND2_X1  g190(.A1(new_n607), .A2(new_n614), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n616), .A2(G868), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n617), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g193(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g194(.A(KEYINPUT3), .B(G2104), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(new_n475), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  INV_X1    g198(.A(G2100), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT79), .Z(new_n626));
  NAND2_X1  g201(.A1(new_n482), .A2(G135), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n484), .A2(G123), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n471), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n627), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  OAI211_X1 g207(.A(new_n626), .B(new_n632), .C1(new_n624), .C2(new_n623), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT80), .Z(G156));
  XNOR2_X1  g209(.A(G2427), .B(G2438), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2430), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT15), .B(G2435), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n638), .A2(KEYINPUT14), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT81), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2451), .B(G2454), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT16), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n641), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  AND3_X1   g224(.A1(new_n648), .A2(new_n649), .A3(G14), .ZN(G401));
  XNOR2_X1  g225(.A(G2084), .B(G2090), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2072), .B(G2078), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n651), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(KEYINPUT17), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n654), .B1(new_n655), .B2(new_n652), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT82), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n652), .A2(new_n653), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n658), .A2(new_n651), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n652), .A2(new_n651), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n657), .B(new_n660), .C1(new_n655), .C2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(new_n624), .ZN(new_n663));
  XOR2_X1   g238(.A(KEYINPUT83), .B(G2096), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(G227));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1956), .B(G2474), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT84), .ZN(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  NAND3_X1  g246(.A1(new_n668), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT20), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n668), .B1(new_n670), .B2(new_n671), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n673), .B(new_n676), .C1(new_n667), .C2(new_n675), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1981), .B(G1986), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT86), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(KEYINPUT85), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n681), .B(new_n684), .ZN(G229));
  AOI22_X1  g260(.A1(new_n482), .A2(G141), .B1(G105), .B2(new_n475), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n484), .A2(G129), .ZN(new_n687));
  NAND3_X1  g262(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n688));
  XOR2_X1   g263(.A(new_n688), .B(KEYINPUT26), .Z(new_n689));
  NAND3_X1  g264(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  OR2_X1    g265(.A1(new_n690), .A2(KEYINPUT92), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(KEYINPUT92), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  OR3_X1    g269(.A1(new_n693), .A2(KEYINPUT93), .A3(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(G29), .A2(G32), .ZN(new_n696));
  OAI211_X1 g271(.A(KEYINPUT93), .B(new_n696), .C1(new_n693), .C2(new_n694), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT27), .B(G1996), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n698), .B(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n694), .A2(G35), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(G162), .B2(new_n694), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT29), .Z(new_n704));
  INV_X1    g279(.A(G2090), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(G34), .ZN(new_n707));
  AOI21_X1  g282(.A(G29), .B1(new_n707), .B2(KEYINPUT24), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(KEYINPUT24), .B2(new_n707), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(new_n479), .B2(new_n694), .ZN(new_n710));
  INV_X1    g285(.A(G2084), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(KEYINPUT91), .B(G1348), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n607), .A2(G16), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(G4), .B2(G16), .ZN(new_n715));
  OAI211_X1 g290(.A(new_n706), .B(new_n712), .C1(new_n713), .C2(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n701), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  AND2_X1   g293(.A1(new_n718), .A2(G5), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G301), .B2(G16), .ZN(new_n720));
  INV_X1    g295(.A(G1961), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n710), .A2(new_n711), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n549), .A2(new_n718), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n718), .A2(G19), .ZN(new_n725));
  OR3_X1    g300(.A1(new_n724), .A2(G1341), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g301(.A(G1341), .B1(new_n724), .B2(new_n725), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n722), .A2(new_n723), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n704), .A2(new_n705), .ZN(new_n729));
  AOI211_X1 g304(.A(new_n728), .B(new_n729), .C1(new_n713), .C2(new_n715), .ZN(new_n730));
  OAI21_X1  g305(.A(KEYINPUT94), .B1(G16), .B2(G21), .ZN(new_n731));
  NOR2_X1   g306(.A1(G286), .A2(new_n718), .ZN(new_n732));
  MUX2_X1   g307(.A(new_n731), .B(KEYINPUT94), .S(new_n732), .Z(new_n733));
  INV_X1    g308(.A(G1966), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n733), .A2(new_n734), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n694), .A2(G26), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n482), .A2(G140), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n484), .A2(G128), .ZN(new_n740));
  OR2_X1    g315(.A1(G104), .A2(G2105), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n741), .B(G2104), .C1(G116), .C2(new_n471), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n738), .B1(new_n744), .B2(new_n694), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2067), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n718), .A2(G20), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT23), .Z(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G299), .B2(G16), .ZN(new_n749));
  INV_X1    g324(.A(G1956), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NOR4_X1   g326(.A1(new_n735), .A2(new_n736), .A3(new_n746), .A4(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n694), .A2(G27), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G164), .B2(new_n694), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(G2078), .ZN(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT30), .B(G28), .ZN(new_n756));
  OR2_X1    g331(.A1(KEYINPUT31), .A2(G11), .ZN(new_n757));
  NAND2_X1  g332(.A1(KEYINPUT31), .A2(G11), .ZN(new_n758));
  AOI22_X1  g333(.A1(new_n756), .A2(new_n694), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n755), .B(new_n759), .C1(new_n694), .C2(new_n631), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n694), .A2(G33), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n762));
  NAND2_X1  g337(.A1(G103), .A2(G2104), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n763), .B2(G2105), .ZN(new_n764));
  NAND4_X1  g339(.A1(new_n471), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n482), .A2(G139), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(G115), .A2(G2104), .ZN(new_n767));
  INV_X1    g342(.A(G127), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n481), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G2105), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n761), .B1(new_n772), .B2(new_n694), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n720), .A2(new_n721), .B1(new_n773), .B2(G2072), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n774), .B1(G2072), .B2(new_n773), .C1(G2078), .C2(new_n754), .ZN(new_n775));
  AOI211_X1 g350(.A(new_n760), .B(new_n775), .C1(new_n750), .C2(new_n749), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n717), .A2(new_n730), .A3(new_n752), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n718), .A2(G22), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n778), .B1(G166), .B2(new_n718), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G1971), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n718), .A2(G23), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G288), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT33), .B(G1976), .ZN(new_n784));
  AND2_X1   g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n781), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n576), .A2(G16), .A3(new_n581), .ZN(new_n788));
  OR2_X1    g363(.A1(G6), .A2(G16), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n790), .A2(KEYINPUT32), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT32), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n788), .A2(new_n792), .A3(new_n789), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n794), .A2(G1981), .ZN(new_n795));
  INV_X1    g370(.A(G1981), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n791), .A2(new_n796), .A3(new_n793), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n779), .A2(G1971), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n787), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n800), .A2(KEYINPUT34), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT34), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n787), .A2(new_n802), .A3(new_n798), .A4(new_n799), .ZN(new_n803));
  XOR2_X1   g378(.A(KEYINPUT35), .B(G1991), .Z(new_n804));
  INV_X1    g379(.A(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n694), .A2(G25), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n482), .A2(G131), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n484), .A2(G119), .ZN(new_n808));
  OR2_X1    g383(.A1(G95), .A2(G2105), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n809), .B(G2104), .C1(G107), .C2(new_n471), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n807), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(KEYINPUT87), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(KEYINPUT87), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n805), .B(new_n806), .C1(new_n814), .C2(new_n694), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n694), .B1(new_n812), .B2(new_n813), .ZN(new_n816));
  INV_X1    g391(.A(new_n806), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n804), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n815), .A2(KEYINPUT88), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(KEYINPUT88), .B1(new_n815), .B2(new_n818), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n718), .A2(G24), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(new_n588), .B2(new_n718), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(G1986), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n820), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n801), .A2(new_n803), .A3(new_n819), .A4(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT89), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n819), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n828), .A2(new_n820), .A3(new_n823), .ZN(new_n829));
  NAND4_X1  g404(.A1(new_n829), .A2(new_n801), .A3(KEYINPUT89), .A4(new_n803), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n827), .A2(KEYINPUT36), .A3(new_n830), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n829), .A2(new_n801), .A3(new_n803), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT36), .ZN(new_n833));
  AOI21_X1  g408(.A(KEYINPUT90), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n777), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n827), .A2(KEYINPUT90), .A3(new_n830), .A4(KEYINPUT36), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(G311));
  NAND2_X1  g412(.A1(new_n831), .A2(new_n834), .ZN(new_n838));
  INV_X1    g413(.A(new_n777), .ZN(new_n839));
  AND4_X1   g414(.A1(KEYINPUT95), .A2(new_n838), .A3(new_n836), .A4(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(KEYINPUT95), .B1(new_n835), .B2(new_n836), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(G150));
  INV_X1    g417(.A(G55), .ZN(new_n843));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  OAI22_X1  g419(.A1(new_n529), .A2(new_n843), .B1(new_n844), .B2(new_n508), .ZN(new_n845));
  AOI22_X1  g420(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(new_n511), .ZN(new_n847));
  OAI21_X1  g422(.A(G860), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT37), .Z(new_n849));
  NOR2_X1   g424(.A1(new_n845), .A2(new_n847), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT96), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(new_n549), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT96), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n850), .B(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n549), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT38), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n857), .B(new_n858), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n606), .A2(new_n614), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n857), .B(KEYINPUT38), .ZN(new_n862));
  INV_X1    g437(.A(new_n860), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n861), .A2(new_n864), .A3(KEYINPUT39), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT97), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT98), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT39), .B1(new_n861), .B2(new_n864), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n869), .A2(G860), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n867), .A2(new_n868), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n868), .B1(new_n867), .B2(new_n870), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n849), .B1(new_n871), .B2(new_n872), .ZN(G145));
  XNOR2_X1  g448(.A(new_n479), .B(new_n488), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(new_n631), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n490), .A2(new_n493), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n498), .A2(KEYINPUT99), .A3(new_n500), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT99), .B1(new_n498), .B2(new_n500), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n876), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AND2_X1   g454(.A1(new_n691), .A2(new_n692), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n744), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n693), .A2(new_n743), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n771), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n771), .B1(new_n881), .B2(new_n882), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI22_X1  g461(.A1(new_n482), .A2(G142), .B1(new_n484), .B2(G130), .ZN(new_n887));
  OAI21_X1  g462(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n888));
  INV_X1    g463(.A(G118), .ZN(new_n889));
  AOI22_X1  g464(.A1(new_n888), .A2(KEYINPUT100), .B1(new_n889), .B2(G2105), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n890), .B1(KEYINPUT100), .B2(new_n888), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n892), .B(new_n622), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n814), .B(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(KEYINPUT101), .B(KEYINPUT102), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n894), .B(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n885), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT99), .ZN(new_n898));
  INV_X1    g473(.A(new_n500), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n499), .B1(new_n620), .B2(new_n496), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n498), .A2(KEYINPUT99), .A3(new_n500), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n494), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n897), .A2(new_n903), .A3(new_n883), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n886), .A2(new_n896), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n886), .A2(new_n904), .ZN(new_n908));
  INV_X1    g483(.A(new_n896), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n905), .A2(new_n906), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n875), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n875), .ZN(new_n914));
  AND2_X1   g489(.A1(new_n905), .A2(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n915), .B2(new_n910), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n913), .A2(KEYINPUT40), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(KEYINPUT40), .B1(new_n913), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(G395));
  XOR2_X1   g494(.A(KEYINPUT105), .B(KEYINPUT42), .Z(new_n920));
  XNOR2_X1  g495(.A(new_n857), .B(new_n616), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n922));
  NAND2_X1  g497(.A1(G299), .A2(new_n606), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(G299), .A2(new_n606), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n921), .A2(new_n922), .A3(new_n926), .ZN(new_n927));
  OR2_X1    g502(.A1(new_n857), .A2(new_n616), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n857), .A2(new_n616), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT41), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n930), .B1(new_n924), .B2(new_n925), .ZN(new_n931));
  INV_X1    g506(.A(new_n925), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n932), .A2(new_n923), .A3(KEYINPUT41), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n928), .A2(new_n929), .A3(new_n931), .A4(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n927), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n922), .B1(new_n921), .B2(new_n926), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n920), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n588), .B(G305), .ZN(new_n938));
  INV_X1    g513(.A(G288), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n939), .A2(G166), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n939), .A2(G166), .ZN(new_n942));
  OR3_X1    g517(.A1(new_n938), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n921), .A2(new_n926), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT104), .ZN(new_n948));
  INV_X1    g523(.A(new_n920), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n948), .A2(new_n949), .A3(new_n934), .A4(new_n927), .ZN(new_n950));
  AND3_X1   g525(.A1(new_n937), .A2(new_n946), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n946), .B1(new_n937), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g527(.A(G868), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n953), .B1(G868), .B2(new_n850), .ZN(G295));
  OAI21_X1  g529(.A(new_n953), .B1(G868), .B2(new_n850), .ZN(G331));
  XNOR2_X1  g530(.A(G301), .B(G168), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n852), .A2(new_n856), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(new_n956), .B1(new_n852), .B2(new_n856), .ZN(new_n959));
  OAI211_X1 g534(.A(new_n931), .B(new_n933), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(new_n959), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n961), .A2(new_n926), .A3(new_n957), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n945), .ZN(new_n964));
  INV_X1    g539(.A(G37), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n960), .A2(new_n946), .A3(new_n962), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n967), .A2(KEYINPUT43), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT43), .ZN(new_n969));
  NAND4_X1  g544(.A1(new_n964), .A2(new_n969), .A3(new_n965), .A4(new_n966), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n972));
  AOI21_X1  g547(.A(KEYINPUT44), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT44), .ZN(new_n974));
  AOI211_X1 g549(.A(KEYINPUT106), .B(new_n974), .C1(new_n968), .C2(new_n970), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n973), .A2(new_n975), .ZN(G397));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n903), .B2(G1384), .ZN(new_n978));
  OAI211_X1 g553(.A(G40), .B(new_n470), .C1(new_n477), .C2(new_n478), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  OR3_X1    g556(.A1(new_n981), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT46), .B1(new_n981), .B2(G1996), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n743), .B(G2067), .ZN(new_n984));
  OR2_X1    g559(.A1(new_n693), .A2(new_n984), .ZN(new_n985));
  AOI22_X1  g560(.A1(new_n982), .A2(new_n983), .B1(new_n980), .B2(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT47), .ZN(new_n987));
  INV_X1    g562(.A(G1996), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n880), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n984), .B1(new_n693), .B2(G1996), .ZN(new_n990));
  AND2_X1   g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n814), .B(new_n805), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n980), .ZN(new_n994));
  XNOR2_X1  g569(.A(new_n994), .B(KEYINPUT126), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n981), .A2(G1986), .A3(G290), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT48), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n991), .A2(new_n804), .A3(new_n814), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(G2067), .B2(new_n743), .ZN(new_n1000));
  AOI211_X1 g575(.A(new_n987), .B(new_n998), .C1(new_n980), .C2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT120), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT50), .ZN(new_n1003));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n879), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n498), .A2(new_n500), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n876), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(new_n1004), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n979), .B1(new_n1008), .B2(KEYINPUT50), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT115), .B(G2084), .ZN(new_n1010));
  AND3_X1   g585(.A1(new_n1005), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1384), .B1(new_n1006), .B2(new_n876), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n979), .B1(KEYINPUT45), .B2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(G1966), .B1(new_n978), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1002), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G168), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT45), .B1(new_n879), .B2(new_n1004), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1012), .A2(KEYINPUT45), .ZN(new_n1019));
  INV_X1    g594(.A(new_n979), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n734), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1005), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1022), .A2(new_n1023), .A3(KEYINPUT120), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1015), .A2(new_n1017), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT51), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1015), .A2(G8), .A3(new_n1024), .ZN(new_n1027));
  XOR2_X1   g602(.A(new_n1017), .B(KEYINPUT121), .Z(new_n1028));
  AOI21_X1  g603(.A(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1016), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n1017), .A2(KEYINPUT51), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(KEYINPUT122), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(G8), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT122), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(new_n1035), .A3(new_n1031), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1025), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT62), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1020), .A2(new_n879), .A3(new_n1004), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n939), .A2(G1976), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1040), .A2(new_n1041), .A3(G8), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(KEYINPUT52), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT110), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT110), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(new_n1045), .A3(KEYINPUT52), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G1976), .ZN(new_n1048));
  AOI21_X1  g623(.A(KEYINPUT52), .B1(G288), .B2(new_n1048), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1040), .A2(new_n1041), .A3(new_n1049), .A4(G8), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n523), .A2(G61), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT73), .ZN(new_n1052));
  XNOR2_X1  g627(.A(new_n577), .B(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n511), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(G1981), .B1(new_n1054), .B2(new_n575), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n522), .A2(G86), .A3(new_n523), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n581), .A2(new_n796), .A3(new_n1056), .A4(new_n573), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1055), .A2(new_n1057), .A3(KEYINPUT111), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT111), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(G1981), .C1(new_n1054), .C2(new_n575), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g636(.A(G8), .B(new_n1040), .C1(new_n1061), .C2(KEYINPUT49), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1061), .A2(KEYINPUT49), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1050), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT108), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT107), .B1(new_n1012), .B2(KEYINPUT45), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT107), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1068), .B(new_n977), .C1(G164), .C2(G1384), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1067), .A2(new_n1020), .A3(new_n1069), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n903), .A2(new_n977), .A3(G1384), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1066), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(G1971), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n977), .B1(G164), .B2(G1384), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n979), .B1(new_n1074), .B2(KEYINPUT107), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n879), .A2(KEYINPUT45), .A3(new_n1004), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(KEYINPUT108), .A3(new_n1076), .A4(new_n1069), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1072), .A2(new_n1073), .A3(new_n1077), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n979), .B1(new_n1003), .B2(new_n1012), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n903), .A2(G1384), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1079), .B1(new_n1080), .B2(new_n1003), .ZN(new_n1081));
  OR2_X1    g656(.A1(new_n1081), .A2(G2090), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1016), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n515), .A2(new_n525), .A3(G8), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT55), .ZN(new_n1085));
  XNOR2_X1  g660(.A(new_n1084), .B(new_n1085), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1047), .B(new_n1065), .C1(new_n1083), .C2(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n1088), .A2(G1961), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  OR4_X1    g665(.A1(new_n1090), .A2(new_n1018), .A3(new_n1021), .A4(G2078), .ZN(new_n1091));
  AOI21_X1  g666(.A(G2078), .B1(new_n1072), .B2(new_n1077), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1089), .B(new_n1091), .C1(new_n1092), .C2(KEYINPUT53), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(G171), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1088), .A2(new_n705), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1078), .A2(new_n1095), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1086), .B(KEYINPUT109), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1096), .A2(G8), .A3(new_n1097), .ZN(new_n1098));
  NOR3_X1   g673(.A1(new_n1087), .A2(new_n1094), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT62), .ZN(new_n1100));
  OAI211_X1 g675(.A(new_n1100), .B(new_n1025), .C1(new_n1029), .C2(new_n1037), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1039), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1086), .B1(new_n1096), .B2(G8), .ZN(new_n1103));
  AOI211_X1 g678(.A(new_n1016), .B(G286), .C1(new_n1022), .C2(new_n1023), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1047), .A2(new_n1065), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(KEYINPUT63), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n939), .A2(new_n1048), .ZN(new_n1107));
  XNOR2_X1  g682(.A(new_n1107), .B(KEYINPUT113), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(new_n1063), .B2(new_n1062), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1057), .B(KEYINPUT112), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT114), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1016), .B1(new_n1080), .B2(new_n1020), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT114), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1109), .A2(new_n1114), .A3(new_n1110), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1112), .A2(new_n1113), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1106), .A2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1047), .A2(new_n1065), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT63), .ZN(new_n1119));
  OAI211_X1 g694(.A(new_n1119), .B(new_n1104), .C1(new_n1083), .C2(new_n1086), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1096), .A2(G8), .A3(new_n1097), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1118), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1117), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1102), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n1125));
  INV_X1    g700(.A(new_n713), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1126), .B1(new_n1005), .B2(new_n1009), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n1040), .A2(G2067), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1127), .A2(new_n1128), .A3(new_n1125), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  XOR2_X1   g707(.A(G299), .B(KEYINPUT57), .Z(new_n1133));
  NAND2_X1  g708(.A1(new_n1081), .A2(new_n750), .ZN(new_n1134));
  XNOR2_X1  g709(.A(KEYINPUT56), .B(G2072), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1075), .A2(new_n1076), .A3(new_n1069), .A4(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1132), .A2(new_n1137), .A3(new_n607), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1133), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT60), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1143), .B(new_n606), .C1(new_n1132), .C2(new_n1144), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT116), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1144), .B1(new_n1147), .B2(new_n1129), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n607), .B1(new_n1148), .B2(KEYINPUT119), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(KEYINPUT119), .ZN(new_n1151));
  AOI22_X1  g726(.A1(new_n1150), .A2(new_n1151), .B1(new_n1144), .B2(new_n1132), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1141), .A2(new_n1137), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT61), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT59), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1075), .A2(new_n988), .A3(new_n1076), .A4(new_n1069), .ZN(new_n1157));
  XOR2_X1   g732(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(G1341), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1040), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n855), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1156), .B1(new_n1161), .B2(KEYINPUT118), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(KEYINPUT118), .ZN(new_n1163));
  XNOR2_X1  g738(.A(new_n1162), .B(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1141), .A2(KEYINPUT61), .A3(new_n1137), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1155), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1142), .B1(new_n1152), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT54), .ZN(new_n1168));
  OAI211_X1 g743(.A(G301), .B(new_n1089), .C1(new_n1092), .C2(KEYINPUT53), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1071), .A2(new_n1090), .A3(G2078), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n979), .A2(KEYINPUT123), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1018), .A2(new_n1171), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n979), .A2(KEYINPUT123), .ZN(new_n1173));
  AOI21_X1  g748(.A(KEYINPUT124), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n979), .A2(KEYINPUT123), .ZN(new_n1175));
  AND4_X1   g750(.A1(KEYINPUT124), .A2(new_n978), .A3(new_n1173), .A4(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1170), .B1(new_n1174), .B2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT125), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  OAI211_X1 g754(.A(KEYINPUT125), .B(new_n1170), .C1(new_n1174), .C2(new_n1176), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1169), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  AND2_X1   g756(.A1(new_n1093), .A2(G171), .ZN(new_n1182));
  OAI21_X1  g757(.A(new_n1168), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  OR2_X1    g758(.A1(new_n1092), .A2(KEYINPUT53), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1184), .A2(G301), .A3(new_n1089), .A4(new_n1091), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1089), .B1(new_n1092), .B2(KEYINPUT53), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1186), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1187));
  OAI211_X1 g762(.A(KEYINPUT54), .B(new_n1185), .C1(new_n1187), .C2(G301), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1087), .A2(new_n1098), .ZN(new_n1189));
  AND4_X1   g764(.A1(new_n1183), .A2(new_n1188), .A3(new_n1038), .A4(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1124), .B1(new_n1167), .B2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(new_n993), .ZN(new_n1192));
  XNOR2_X1  g767(.A(new_n588), .B(G1986), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n981), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1001), .B1(new_n1191), .B2(new_n1194), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g770(.A1(new_n913), .A2(new_n916), .ZN(new_n1197));
  NOR2_X1   g771(.A1(G229), .A2(G401), .ZN(new_n1198));
  NOR2_X1   g772(.A1(G227), .A2(new_n457), .ZN(new_n1199));
  XNOR2_X1  g773(.A(new_n1199), .B(KEYINPUT127), .ZN(new_n1200));
  AND4_X1   g774(.A1(new_n1197), .A2(new_n1198), .A3(new_n1200), .A4(new_n971), .ZN(G308));
  NAND4_X1  g775(.A1(new_n1197), .A2(new_n1198), .A3(new_n1200), .A4(new_n971), .ZN(G225));
endmodule


