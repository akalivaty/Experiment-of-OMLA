//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:38 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009;
  NOR2_X1   g000(.A1(G475), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G125), .ZN(new_n188));
  NOR3_X1   g002(.A1(new_n188), .A2(KEYINPUT16), .A3(G140), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(G125), .A2(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n196));
  OAI211_X1 g010(.A(G146), .B(new_n190), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n196), .B1(new_n192), .B2(new_n193), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n198), .B1(new_n199), .B2(new_n189), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT74), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n197), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  OAI211_X1 g016(.A(KEYINPUT74), .B(new_n198), .C1(new_n199), .C2(new_n189), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(G237), .A2(G953), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(G143), .A3(G214), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(G143), .B1(new_n205), .B2(G214), .ZN(new_n208));
  OAI21_X1  g022(.A(G131), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n205), .A2(G214), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G131), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(new_n206), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n209), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  OR2_X1    g030(.A1(new_n209), .A2(new_n215), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n204), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G113), .B(G122), .ZN(new_n219));
  INV_X1    g033(.A(G104), .ZN(new_n220));
  XNOR2_X1  g034(.A(new_n219), .B(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n194), .A2(KEYINPUT76), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT76), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n192), .A2(new_n223), .A3(new_n193), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n222), .A2(new_n198), .A3(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n195), .A2(G146), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT18), .A2(G131), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n228), .B1(new_n207), .B2(new_n208), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n212), .A2(KEYINPUT18), .A3(G131), .A4(new_n206), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n227), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n218), .A2(new_n221), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n199), .A2(new_n189), .ZN(new_n234));
  AOI22_X1  g048(.A1(new_n209), .A2(new_n214), .B1(new_n234), .B2(G146), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT91), .ZN(new_n236));
  AOI21_X1  g050(.A(KEYINPUT19), .B1(new_n224), .B2(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(KEYINPUT76), .B1(new_n236), .B2(KEYINPUT19), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(new_n192), .B2(new_n193), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n198), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n235), .A2(new_n240), .B1(new_n227), .B2(new_n231), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT92), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n221), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n244), .B1(new_n241), .B2(KEYINPUT92), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n233), .B(KEYINPUT93), .C1(new_n243), .C2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n235), .A2(new_n240), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n232), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT92), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n242), .A3(new_n244), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT93), .B1(new_n252), .B2(new_n233), .ZN(new_n253));
  OAI211_X1 g067(.A(KEYINPUT20), .B(new_n187), .C1(new_n247), .C2(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n233), .B1(new_n243), .B2(new_n245), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(new_n187), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT20), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n218), .A2(new_n232), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n244), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(new_n233), .ZN(new_n261));
  INV_X1    g075(.A(G902), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G475), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n254), .A2(new_n258), .A3(new_n264), .ZN(new_n265));
  XOR2_X1   g079(.A(KEYINPUT9), .B(G234), .Z(new_n266));
  INV_X1    g080(.A(G953), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(G217), .A3(new_n267), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n268), .B(KEYINPUT95), .Z(new_n269));
  XNOR2_X1  g083(.A(G128), .B(G143), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT13), .ZN(new_n271));
  INV_X1    g085(.A(G128), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n272), .A2(KEYINPUT13), .A3(G143), .ZN(new_n273));
  INV_X1    g087(.A(G134), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n271), .A2(new_n275), .B1(new_n274), .B2(new_n270), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT94), .ZN(new_n277));
  INV_X1    g091(.A(G122), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n277), .B1(new_n278), .B2(G116), .ZN(new_n279));
  INV_X1    g093(.A(G116), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT94), .A3(G122), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n279), .A2(new_n281), .B1(G116), .B2(new_n278), .ZN(new_n282));
  INV_X1    g096(.A(G107), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n282), .A2(new_n283), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n276), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n278), .A2(G116), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n283), .B1(new_n287), .B2(KEYINPUT14), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n282), .B(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(new_n270), .B(new_n274), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n269), .A2(new_n286), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n269), .B1(new_n286), .B2(new_n291), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G478), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n295), .B(new_n262), .C1(KEYINPUT15), .C2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n294), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(new_n262), .A3(new_n292), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n296), .A2(KEYINPUT15), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G952), .ZN(new_n304));
  AOI211_X1 g118(.A(G953), .B(new_n304), .C1(G234), .C2(G237), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n262), .B(new_n267), .C1(G234), .C2(G237), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT21), .B(G898), .Z(new_n309));
  OAI21_X1  g123(.A(new_n306), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  XOR2_X1   g124(.A(new_n310), .B(KEYINPUT96), .Z(new_n311));
  NAND2_X1  g125(.A1(new_n303), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT97), .B1(new_n265), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n187), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT93), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n255), .A2(new_n315), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n314), .B1(new_n316), .B2(new_n246), .ZN(new_n317));
  AOI22_X1  g131(.A1(new_n317), .A2(KEYINPUT20), .B1(G475), .B2(new_n263), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT97), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n297), .A2(new_n301), .A3(new_n311), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n318), .A2(new_n319), .A3(new_n258), .A4(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n313), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(G214), .B1(G237), .B2(G902), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT2), .ZN(new_n325));
  INV_X1    g139(.A(G113), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(new_n326), .A3(KEYINPUT65), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT65), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(KEYINPUT2), .B2(G113), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n327), .A2(new_n329), .B1(KEYINPUT2), .B2(G113), .ZN(new_n330));
  XNOR2_X1  g144(.A(G116), .B(G119), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n330), .B(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT3), .B1(new_n220), .B2(G107), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT3), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(new_n283), .A3(G104), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n220), .A2(G107), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(KEYINPUT82), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT82), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n334), .A2(new_n336), .A3(new_n340), .A4(new_n337), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(G101), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G101), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n334), .A2(new_n336), .A3(new_n343), .A4(new_n337), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT4), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND4_X1  g160(.A1(new_n339), .A2(KEYINPUT4), .A3(G101), .A4(new_n341), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n333), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G119), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G116), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n280), .A2(G119), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n350), .A2(new_n351), .A3(KEYINPUT5), .ZN(new_n352));
  OAI21_X1  g166(.A(G113), .B1(new_n350), .B2(KEYINPUT5), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT85), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n331), .A2(KEYINPUT5), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n280), .A2(G119), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT5), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n326), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n355), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n330), .A2(new_n331), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n354), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n337), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n220), .A2(G107), .ZN(new_n364));
  OAI21_X1  g178(.A(G101), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n344), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n348), .A2(new_n367), .ZN(new_n368));
  XOR2_X1   g182(.A(G110), .B(G122), .Z(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n369), .B1(new_n348), .B2(new_n367), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(KEYINPUT6), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n198), .A2(G143), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n211), .A2(G146), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT0), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(new_n272), .ZN(new_n378));
  NOR2_X1   g192(.A1(KEYINPUT0), .A2(G128), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n376), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(G143), .B(G146), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n381), .B1(new_n377), .B2(new_n272), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n188), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n374), .A2(G128), .ZN(new_n384));
  INV_X1    g198(.A(new_n384), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n272), .A2(KEYINPUT1), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(new_n375), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(KEYINPUT64), .B1(new_n381), .B2(new_n386), .ZN(new_n389));
  AND4_X1   g203(.A1(KEYINPUT64), .A2(new_n386), .A3(new_n374), .A4(new_n375), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n385), .B(new_n388), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n383), .B1(new_n391), .B2(new_n188), .ZN(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT87), .B(G224), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n267), .ZN(new_n394));
  XOR2_X1   g208(.A(new_n392), .B(new_n394), .Z(new_n395));
  INV_X1    g209(.A(KEYINPUT6), .ZN(new_n396));
  OAI211_X1 g210(.A(new_n396), .B(new_n369), .C1(new_n348), .C2(new_n367), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n397), .A2(new_n398), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n373), .B(new_n395), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n392), .B1(KEYINPUT89), .B2(KEYINPUT7), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n394), .A2(KEYINPUT7), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  OR2_X1    g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n355), .B(KEYINPUT88), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n361), .B1(new_n406), .B2(new_n353), .ZN(new_n407));
  INV_X1    g221(.A(new_n366), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n369), .B(KEYINPUT8), .Z(new_n410));
  OAI211_X1 g224(.A(new_n409), .B(new_n410), .C1(new_n408), .C2(new_n362), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n402), .A2(new_n404), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n405), .A2(new_n371), .A3(new_n411), .A4(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n401), .A2(new_n262), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT90), .ZN(new_n415));
  OAI21_X1  g229(.A(G210), .B1(G237), .B2(G902), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n348), .A2(new_n367), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n419), .A2(KEYINPUT86), .A3(new_n396), .A4(new_n369), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n397), .A2(new_n398), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n396), .B1(new_n368), .B2(new_n370), .ZN(new_n422));
  AOI22_X1  g236(.A1(new_n420), .A2(new_n421), .B1(new_n422), .B2(new_n372), .ZN(new_n423));
  AOI21_X1  g237(.A(G902), .B1(new_n423), .B2(new_n395), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n417), .A2(new_n415), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n413), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n324), .B1(new_n418), .B2(new_n426), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n322), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(KEYINPUT78), .B(KEYINPUT79), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n430));
  XNOR2_X1  g244(.A(new_n429), .B(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT22), .B(G137), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT72), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n434), .B1(new_n349), .B2(G128), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n349), .A2(G128), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(KEYINPUT23), .A3(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT23), .B1(new_n272), .B2(G119), .ZN(new_n438));
  AOI21_X1  g252(.A(KEYINPUT72), .B1(new_n272), .B2(G119), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G110), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n437), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT75), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(KEYINPUT24), .A2(G110), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(KEYINPUT24), .A2(G110), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(KEYINPUT71), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT71), .ZN(new_n449));
  INV_X1    g263(.A(new_n447), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n449), .B1(new_n450), .B2(new_n445), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT70), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n453), .B1(new_n349), .B2(G128), .ZN(new_n454));
  NOR3_X1   g268(.A1(new_n272), .A2(KEYINPUT70), .A3(G119), .ZN(new_n455));
  OAI22_X1  g269(.A1(new_n454), .A2(new_n455), .B1(new_n349), .B2(G128), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n437), .A2(new_n440), .A3(KEYINPUT75), .A4(new_n441), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n444), .A2(new_n457), .A3(new_n458), .ZN(new_n459));
  AND2_X1   g273(.A1(new_n197), .A2(new_n225), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT77), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT77), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n437), .A2(new_n440), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT73), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n437), .A2(new_n440), .A3(KEYINPUT73), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(G110), .A3(new_n469), .ZN(new_n470));
  OR2_X1    g284(.A1(new_n452), .A2(new_n456), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n470), .A2(new_n202), .A3(new_n471), .A4(new_n203), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n433), .B1(new_n465), .B2(new_n472), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n459), .A2(new_n460), .A3(KEYINPUT77), .ZN(new_n474));
  AOI21_X1  g288(.A(KEYINPUT77), .B1(new_n459), .B2(new_n460), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n472), .B(new_n433), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT80), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT25), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n479), .A2(new_n480), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n478), .A2(new_n262), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n485));
  INV_X1    g299(.A(new_n433), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n476), .ZN(new_n488));
  OAI211_X1 g302(.A(KEYINPUT80), .B(KEYINPUT25), .C1(new_n488), .C2(G902), .ZN(new_n489));
  INV_X1    g303(.A(G217), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(G234), .B2(new_n262), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n484), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT81), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n484), .A2(new_n489), .A3(KEYINPUT81), .A4(new_n491), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n491), .A2(G902), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n478), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n499), .B(G101), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n205), .A2(G210), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n274), .A2(G137), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n274), .A2(G137), .ZN(new_n505));
  OAI21_X1  g319(.A(G131), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT11), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n274), .B2(G137), .ZN(new_n508));
  INV_X1    g322(.A(G137), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(KEYINPUT11), .A3(G134), .ZN(new_n510));
  NAND4_X1  g324(.A1(new_n508), .A2(new_n510), .A3(new_n213), .A4(new_n503), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n508), .A2(new_n503), .A3(new_n510), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(G131), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n511), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n380), .A2(new_n382), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n391), .A2(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n333), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT67), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n516), .A2(new_n517), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n386), .A2(new_n374), .A3(new_n375), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT64), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n386), .A2(new_n374), .A3(new_n375), .A4(KEYINPUT64), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n384), .B(new_n387), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n521), .B1(new_n526), .B2(new_n512), .ZN(new_n527));
  INV_X1    g341(.A(new_n333), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n520), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR3_X1   g343(.A1(new_n518), .A2(KEYINPUT67), .A3(new_n333), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n519), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(KEYINPUT28), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n527), .A2(new_n528), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n533), .A2(KEYINPUT28), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n502), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n387), .B1(new_n524), .B2(new_n525), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n512), .B1(new_n537), .B2(new_n385), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n515), .A2(new_n511), .B1(new_n380), .B2(new_n382), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT30), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n391), .A2(new_n513), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT30), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n542), .A3(new_n521), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n540), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n533), .B1(new_n544), .B2(new_n528), .ZN(new_n545));
  AOI21_X1  g359(.A(KEYINPUT66), .B1(new_n545), .B2(new_n502), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n333), .B1(new_n540), .B2(new_n543), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT66), .ZN(new_n548));
  INV_X1    g362(.A(new_n502), .ZN(new_n549));
  NOR4_X1   g363(.A1(new_n547), .A2(new_n548), .A3(new_n533), .A4(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT31), .ZN(new_n551));
  NOR3_X1   g365(.A1(new_n546), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NOR3_X1   g366(.A1(new_n538), .A2(KEYINPUT30), .A3(new_n539), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n542), .B1(new_n541), .B2(new_n521), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n528), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n555), .A2(new_n519), .A3(new_n502), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n551), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n536), .B1(new_n552), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT32), .ZN(new_n560));
  INV_X1    g374(.A(G472), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(new_n262), .A3(KEYINPUT68), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT68), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(G472), .B2(G902), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n559), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n556), .A2(new_n548), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n545), .A2(KEYINPUT66), .A3(new_n502), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n567), .A2(KEYINPUT31), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n535), .B1(new_n569), .B2(new_n557), .ZN(new_n570));
  INV_X1    g384(.A(new_n565), .ZN(new_n571));
  OAI21_X1  g385(.A(KEYINPUT32), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n532), .A2(new_n534), .A3(new_n502), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT29), .ZN(new_n575));
  INV_X1    g389(.A(new_n545), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n549), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n574), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n527), .A2(new_n528), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n519), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT28), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT69), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT69), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n583), .A3(KEYINPUT28), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n582), .A2(KEYINPUT29), .A3(new_n534), .A4(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n262), .B1(new_n585), .B2(new_n549), .ZN(new_n586));
  OAI21_X1  g400(.A(G472), .B1(new_n578), .B2(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n498), .B1(new_n573), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(G221), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n266), .B2(new_n262), .ZN(new_n590));
  XNOR2_X1  g404(.A(G110), .B(G140), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n267), .A2(G227), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n591), .B(new_n592), .Z(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT10), .B1(new_n526), .B2(new_n366), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n391), .A2(new_n596), .A3(new_n408), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n516), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n346), .A2(new_n347), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n517), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n599), .B1(new_n598), .B2(new_n601), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n594), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(KEYINPUT83), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT83), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n606), .B(new_n594), .C1(new_n602), .C2(new_n603), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n526), .A2(new_n366), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n391), .A2(new_n408), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n516), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT12), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n602), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n612), .A2(new_n613), .A3(new_n593), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n605), .A2(new_n607), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(G469), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n262), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT84), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT84), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n615), .A2(new_n619), .A3(new_n616), .A4(new_n262), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  OR3_X1    g435(.A1(new_n602), .A2(new_n603), .A3(new_n594), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n612), .A2(new_n613), .ZN(new_n623));
  OAI211_X1 g437(.A(G469), .B(new_n622), .C1(new_n623), .C2(new_n593), .ZN(new_n624));
  NAND2_X1  g438(.A1(G469), .A2(G902), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n590), .B1(new_n621), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n428), .A2(new_n588), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(KEYINPUT98), .B(G101), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT99), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n629), .B(new_n631), .ZN(G3));
  INV_X1    g446(.A(new_n498), .ZN(new_n633));
  OAI21_X1  g447(.A(G472), .B1(new_n570), .B2(G902), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n559), .A2(new_n565), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n628), .A2(new_n633), .A3(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n295), .A2(KEYINPUT33), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT33), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n293), .A2(new_n294), .A3(new_n640), .ZN(new_n641));
  OAI211_X1 g455(.A(G478), .B(new_n262), .C1(new_n639), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n299), .A2(new_n296), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n265), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n416), .A2(KEYINPUT100), .ZN(new_n646));
  OR2_X1    g460(.A1(new_n416), .A2(KEYINPUT100), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n424), .A2(new_n413), .A3(new_n646), .A4(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n414), .A2(KEYINPUT100), .A3(new_n416), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n648), .A2(new_n649), .A3(new_n323), .A4(new_n311), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n638), .A2(new_n645), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT34), .B(G104), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G6));
  INV_X1    g467(.A(new_n317), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(new_n257), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n318), .A3(new_n302), .ZN(new_n656));
  NOR3_X1   g470(.A1(new_n650), .A2(KEYINPUT101), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g472(.A(KEYINPUT101), .B1(new_n650), .B2(new_n656), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n638), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT35), .B(G107), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G9));
  NOR2_X1   g476(.A1(new_n486), .A2(KEYINPUT36), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n485), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(new_n496), .ZN(new_n665));
  AND3_X1   g479(.A1(new_n494), .A2(new_n495), .A3(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n636), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n428), .A2(new_n667), .A3(new_n628), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT37), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(new_n441), .ZN(G12));
  NAND3_X1  g484(.A1(new_n648), .A2(new_n649), .A3(new_n323), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n671), .B1(new_n573), .B2(new_n587), .ZN(new_n672));
  INV_X1    g486(.A(new_n666), .ZN(new_n673));
  OR2_X1    g487(.A1(new_n308), .A2(G900), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n306), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n656), .A2(new_n676), .ZN(new_n677));
  AND4_X1   g491(.A1(new_n628), .A2(new_n672), .A3(new_n673), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(new_n272), .ZN(G30));
  XNOR2_X1  g493(.A(new_n675), .B(KEYINPUT39), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n628), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n681), .A2(KEYINPUT40), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n418), .A2(new_n426), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT38), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n265), .A2(new_n302), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n666), .A2(new_n690), .A3(new_n323), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n687), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  OR2_X1    g506(.A1(new_n691), .A2(new_n688), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n546), .A2(new_n550), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n580), .A2(new_n549), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(KEYINPUT102), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n561), .B1(new_n698), .B2(new_n262), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n573), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n692), .A2(new_n693), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT104), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n692), .A2(new_n693), .A3(KEYINPUT104), .A4(new_n701), .ZN(new_n705));
  AOI211_X1 g519(.A(new_n683), .B(new_n684), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n211), .ZN(G45));
  NOR2_X1   g521(.A1(new_n645), .A2(new_n676), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n672), .A2(new_n628), .A3(new_n673), .A4(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n626), .B1(new_n618), .B2(new_n620), .ZN(new_n712));
  NOR3_X1   g526(.A1(new_n712), .A2(new_n666), .A3(new_n590), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n713), .A2(KEYINPUT105), .A3(new_n672), .A4(new_n708), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  AOI21_X1  g530(.A(new_n616), .B1(new_n615), .B2(new_n262), .ZN(new_n717));
  AOI211_X1 g531(.A(new_n590), .B(new_n717), .C1(new_n618), .C2(new_n620), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n573), .A2(new_n587), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n650), .A2(new_n645), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n718), .A2(new_n719), .A3(new_n633), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT41), .B(G113), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G15));
  INV_X1    g537(.A(new_n659), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n588), .B(new_n718), .C1(new_n724), .C2(new_n657), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  AND3_X1   g540(.A1(new_n648), .A2(new_n649), .A3(new_n323), .ZN(new_n727));
  INV_X1    g541(.A(new_n590), .ZN(new_n728));
  INV_X1    g542(.A(new_n717), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n727), .A2(new_n621), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT106), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n717), .B1(new_n618), .B2(new_n620), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n733), .A2(KEYINPUT106), .A3(new_n728), .A4(new_n727), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n666), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n719), .A2(new_n322), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  AND3_X1   g552(.A1(new_n582), .A2(new_n534), .A3(new_n584), .ZN(new_n739));
  OAI22_X1  g553(.A1(new_n552), .A2(new_n558), .B1(new_n739), .B2(new_n502), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n565), .B(KEYINPUT107), .Z(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n634), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n743), .A2(new_n498), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n650), .A2(new_n689), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n744), .A2(new_n718), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  INV_X1    g561(.A(new_n708), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n743), .ZN(new_n749));
  AOI21_X1  g563(.A(KEYINPUT106), .B1(new_n718), .B2(new_n727), .ZN(new_n750));
  INV_X1    g564(.A(new_n734), .ZN(new_n751));
  OAI211_X1 g565(.A(new_n673), .B(new_n749), .C1(new_n750), .C2(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT108), .B(G125), .Z(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G27));
  INV_X1    g568(.A(new_n624), .ZN(new_n755));
  XOR2_X1   g569(.A(new_n625), .B(KEYINPUT109), .Z(new_n756));
  AOI211_X1 g570(.A(new_n755), .B(new_n756), .C1(new_n618), .C2(new_n620), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n590), .A2(new_n324), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n418), .A2(new_n426), .A3(new_n759), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n757), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n756), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n621), .A2(new_n624), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n760), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT110), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n588), .B(new_n708), .C1(new_n761), .C2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(KEYINPUT111), .A2(KEYINPUT42), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n588), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n758), .B1(new_n757), .B2(new_n760), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n763), .A2(new_n764), .A3(KEYINPUT110), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n767), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n772), .A2(new_n708), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G131), .ZN(G33));
  NAND2_X1  g590(.A1(new_n772), .A2(new_n677), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  NOR2_X1   g592(.A1(new_n685), .A2(new_n324), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n642), .A2(new_n643), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n265), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(KEYINPUT43), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(new_n636), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(KEYINPUT44), .A3(new_n673), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n784), .A2(KEYINPUT112), .A3(KEYINPUT44), .A4(new_n673), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n780), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT44), .B1(new_n784), .B2(new_n673), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n622), .B1(new_n623), .B2(new_n593), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n793), .A2(G469), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n762), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT46), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n795), .A2(KEYINPUT46), .A3(new_n762), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n798), .A2(new_n621), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n800), .A2(new_n728), .A3(new_n680), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n790), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n789), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  NAND2_X1  g618(.A1(new_n800), .A2(new_n728), .ZN(new_n805));
  XOR2_X1   g619(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(KEYINPUT113), .A2(KEYINPUT47), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n800), .B2(new_n728), .ZN(new_n809));
  NOR3_X1   g623(.A1(new_n807), .A2(new_n748), .A3(new_n809), .ZN(new_n810));
  NOR3_X1   g624(.A1(new_n719), .A2(new_n780), .A3(new_n633), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  INV_X1    g627(.A(new_n678), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n763), .A2(new_n701), .A3(new_n666), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n671), .A2(new_n689), .ZN(new_n816));
  XOR2_X1   g630(.A(new_n675), .B(KEYINPUT115), .Z(new_n817));
  NAND4_X1  g631(.A1(new_n815), .A2(new_n728), .A3(new_n816), .A4(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n715), .A2(new_n814), .A3(new_n752), .A4(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT52), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n678), .B1(new_n711), .B2(new_n714), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(KEYINPUT52), .A3(new_n752), .A4(new_n818), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT116), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n766), .A2(new_n767), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n773), .B1(new_n772), .B2(new_n708), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n777), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n721), .A2(new_n746), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n735), .B2(new_n736), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n628), .B(new_n428), .C1(new_n588), .C2(new_n667), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n645), .B1(new_n265), .B2(new_n303), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n834), .A2(new_n427), .A3(new_n311), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(new_n628), .A3(new_n633), .A4(new_n637), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n833), .A2(KEYINPUT114), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT114), .B1(new_n833), .B2(new_n836), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n832), .B(new_n725), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n749), .B1(new_n761), .B2(new_n765), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n676), .B(new_n760), .C1(new_n573), .C2(new_n587), .ZN(new_n841));
  INV_X1    g655(.A(new_n712), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n655), .A2(new_n318), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n841), .A2(new_n842), .A3(new_n303), .A4(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n666), .B1(new_n840), .B2(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n830), .A2(new_n839), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n821), .A2(new_n823), .A3(KEYINPUT116), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n826), .A2(new_n827), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n824), .ZN(new_n849));
  INV_X1    g663(.A(new_n725), .ZN(new_n850));
  INV_X1    g664(.A(new_n838), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n833), .A2(KEYINPUT114), .A3(new_n836), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n768), .A2(new_n774), .B1(new_n677), .B2(new_n772), .ZN(new_n854));
  INV_X1    g668(.A(new_n845), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n853), .A2(new_n854), .A3(new_n855), .A4(new_n832), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT53), .B1(new_n849), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n848), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT54), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n783), .A2(new_n305), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT117), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n718), .A2(new_n779), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n862), .A2(new_n588), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n864), .B(KEYINPUT48), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n304), .A2(G953), .ZN(new_n866));
  AND2_X1   g680(.A1(new_n862), .A2(new_n744), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n732), .A2(new_n734), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT119), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n867), .A2(KEYINPUT119), .A3(new_n868), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n865), .B(new_n866), .C1(new_n869), .C2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(new_n743), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n862), .A2(new_n673), .A3(new_n872), .A4(new_n863), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT118), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n733), .A2(new_n590), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n876), .B1(new_n807), .B2(new_n809), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n877), .A2(new_n779), .A3(new_n867), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n701), .A2(new_n498), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n863), .A2(new_n305), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n881), .A2(new_n258), .A3(new_n318), .A4(new_n781), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT51), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n687), .A2(new_n718), .A3(new_n744), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n862), .A2(new_n324), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT50), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n862), .A2(new_n886), .A3(KEYINPUT50), .A4(new_n324), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n875), .A2(new_n883), .A3(new_n884), .A4(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n891), .A2(new_n878), .A3(new_n882), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT51), .B1(new_n893), .B2(new_n874), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n871), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n846), .A2(new_n827), .A3(new_n824), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n821), .A2(KEYINPUT116), .A3(new_n823), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT116), .B1(new_n821), .B2(new_n823), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n898), .A3(new_n856), .ZN(new_n899));
  OAI211_X1 g713(.A(KEYINPUT54), .B(new_n896), .C1(new_n899), .C2(new_n827), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n860), .A2(new_n895), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n880), .A2(new_n645), .ZN(new_n902));
  OAI22_X1  g716(.A1(new_n901), .A2(new_n902), .B1(G952), .B2(G953), .ZN(new_n903));
  INV_X1    g717(.A(new_n687), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT49), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n733), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n904), .A2(new_n701), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n733), .A2(new_n905), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n907), .A2(new_n759), .A3(new_n782), .A4(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n903), .B1(new_n498), .B2(new_n909), .ZN(G75));
  XOR2_X1   g724(.A(new_n423), .B(KEYINPUT120), .Z(new_n911));
  XNOR2_X1  g725(.A(KEYINPUT121), .B(KEYINPUT55), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n395), .B(new_n912), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n911), .B(new_n913), .Z(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n848), .A2(new_n857), .A3(G210), .A4(G902), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n915), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n304), .A2(G953), .ZN(new_n919));
  XOR2_X1   g733(.A(new_n919), .B(KEYINPUT123), .Z(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n916), .A2(KEYINPUT122), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(KEYINPUT56), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n914), .B1(new_n916), .B2(KEYINPUT122), .ZN(new_n924));
  AOI211_X1 g738(.A(new_n918), .B(new_n921), .C1(new_n923), .C2(new_n924), .ZN(G51));
  XNOR2_X1  g739(.A(new_n756), .B(KEYINPUT57), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n848), .A2(KEYINPUT54), .A3(new_n857), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT54), .B1(new_n848), .B2(new_n857), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n926), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n615), .ZN(new_n930));
  OR3_X1    g744(.A1(new_n858), .A2(new_n262), .A3(new_n795), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n921), .B1(new_n930), .B2(new_n931), .ZN(G54));
  NOR2_X1   g746(.A1(new_n858), .A2(new_n262), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n933), .A2(KEYINPUT58), .A3(G475), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n316), .A2(new_n246), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(new_n935), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n933), .A2(KEYINPUT58), .A3(G475), .A4(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n921), .B1(new_n936), .B2(new_n938), .ZN(G60));
  NOR2_X1   g753(.A1(new_n639), .A2(new_n641), .ZN(new_n940));
  NAND2_X1  g754(.A1(G478), .A2(G902), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT59), .Z(new_n942));
  NOR2_X1   g756(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(new_n927), .B2(new_n928), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI211_X1 g760(.A(KEYINPUT124), .B(new_n943), .C1(new_n927), .C2(new_n928), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n942), .B1(new_n860), .B2(new_n900), .ZN(new_n949));
  INV_X1    g763(.A(new_n940), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n920), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n948), .A2(new_n951), .ZN(G63));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT60), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n848), .A2(new_n857), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n488), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n848), .A2(new_n857), .A3(new_n664), .A4(new_n955), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n957), .A2(new_n920), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(KEYINPUT61), .B1(new_n958), .B2(KEYINPUT125), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(G66));
  AOI21_X1  g775(.A(new_n267), .B1(new_n309), .B2(new_n393), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n962), .B1(new_n839), .B2(new_n267), .ZN(new_n963));
  INV_X1    g777(.A(G898), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n911), .B1(new_n964), .B2(G953), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n963), .B(new_n965), .ZN(G69));
  INV_X1    g780(.A(KEYINPUT127), .ZN(new_n967));
  AOI22_X1  g781(.A1(new_n810), .A2(new_n811), .B1(new_n789), .B2(new_n802), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n822), .A2(new_n752), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n801), .A2(new_n769), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n969), .B1(new_n970), .B2(new_n816), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n968), .A2(new_n267), .A3(new_n854), .A4(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n237), .A2(new_n239), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n544), .B(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(G900), .A2(G953), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n972), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n684), .B1(new_n704), .B2(new_n705), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n682), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT62), .ZN(new_n980));
  NAND4_X1  g794(.A1(new_n979), .A2(new_n980), .A3(new_n752), .A4(new_n822), .ZN(new_n981));
  OAI21_X1  g795(.A(KEYINPUT62), .B1(new_n706), .B2(new_n969), .ZN(new_n982));
  INV_X1    g796(.A(new_n681), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n983), .A2(new_n588), .A3(new_n779), .A4(new_n834), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n981), .A2(new_n982), .A3(new_n984), .A4(new_n968), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n985), .A2(new_n267), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n977), .B1(new_n986), .B2(new_n975), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n267), .B1(G227), .B2(G900), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n967), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n975), .B1(new_n985), .B2(new_n267), .ZN(new_n990));
  INV_X1    g804(.A(new_n977), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n967), .B(new_n988), .C1(new_n990), .C2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n990), .A2(new_n991), .ZN(new_n994));
  INV_X1    g808(.A(new_n988), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT126), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT126), .ZN(new_n997));
  NOR4_X1   g811(.A1(new_n990), .A2(new_n991), .A3(new_n997), .A4(new_n988), .ZN(new_n998));
  OAI22_X1  g812(.A1(new_n989), .A2(new_n993), .B1(new_n996), .B2(new_n998), .ZN(G72));
  OR2_X1    g813(.A1(new_n899), .A2(new_n827), .ZN(new_n1000));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT63), .Z(new_n1002));
  NAND2_X1  g816(.A1(new_n695), .A2(new_n577), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n1000), .A2(new_n896), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n1002), .B1(new_n985), .B2(new_n839), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1005), .A2(new_n502), .A3(new_n576), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n968), .A2(new_n854), .A3(new_n971), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1002), .B1(new_n1007), .B2(new_n839), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n1008), .A2(new_n549), .A3(new_n545), .ZN(new_n1009));
  AND4_X1   g823(.A1(new_n920), .A2(new_n1004), .A3(new_n1006), .A4(new_n1009), .ZN(G57));
endmodule


