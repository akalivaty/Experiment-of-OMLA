//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n830, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1061, new_n1062, new_n1063, new_n1064, new_n1065, new_n1066,
    new_n1067, new_n1068, new_n1070, new_n1071, new_n1072, new_n1073,
    new_n1074, new_n1075, new_n1076, new_n1077, new_n1078, new_n1079,
    new_n1080, new_n1081, new_n1082, new_n1083, new_n1084;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G104), .ZN(new_n193));
  INV_X1    g007(.A(G101), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n189), .A2(G107), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n190), .A2(new_n193), .A3(new_n194), .A4(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n189), .A2(G107), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n192), .A2(G104), .ZN(new_n198));
  OAI21_X1  g012(.A(G101), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n196), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT77), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT77), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n196), .A2(new_n199), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G113), .ZN(new_n204));
  INV_X1    g018(.A(G116), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G119), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT5), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G116), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(G119), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n211), .A3(KEYINPUT5), .ZN(new_n212));
  XNOR2_X1  g026(.A(G116), .B(G119), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n204), .A2(KEYINPUT2), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(G113), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n208), .A2(new_n212), .B1(new_n213), .B2(new_n217), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n201), .A2(new_n203), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n190), .A2(new_n193), .A3(new_n195), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT74), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT4), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n190), .A2(new_n193), .A3(KEYINPUT74), .A4(new_n195), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n222), .A2(new_n223), .A3(G101), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n210), .A2(new_n211), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(new_n214), .A3(new_n216), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n217), .A2(new_n213), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n196), .A2(KEYINPUT4), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n194), .B1(new_n220), .B2(new_n221), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n231), .B1(new_n232), .B2(new_n224), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n219), .B1(new_n230), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G110), .B(G122), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n235), .B(new_n219), .C1(new_n230), .C2(new_n233), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(KEYINPUT6), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G224), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(G953), .ZN(new_n241));
  INV_X1    g055(.A(G146), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G143), .ZN(new_n243));
  INV_X1    g057(.A(G143), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G146), .ZN(new_n245));
  AOI21_X1  g059(.A(G128), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n244), .A2(KEYINPUT1), .A3(G146), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G128), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(KEYINPUT1), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(new_n243), .A3(new_n245), .ZN(new_n252));
  AOI21_X1  g066(.A(G125), .B1(new_n249), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G125), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n243), .A2(new_n245), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT0), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(new_n250), .ZN(new_n257));
  NOR2_X1   g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G143), .B(G146), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n260), .B1(new_n256), .B2(new_n250), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n254), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n241), .B1(new_n253), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n259), .A2(new_n261), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G125), .ZN(new_n265));
  INV_X1    g079(.A(new_n241), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n252), .B(new_n247), .C1(G128), .C2(new_n260), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n254), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT6), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n234), .A2(new_n271), .A3(new_n236), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n239), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n200), .ZN(new_n274));
  OAI21_X1  g088(.A(KEYINPUT79), .B1(new_n274), .B2(new_n218), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n208), .A2(new_n212), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n228), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT79), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n277), .A2(new_n278), .A3(new_n200), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n219), .A2(new_n275), .A3(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n235), .B(KEYINPUT8), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT7), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n265), .A2(new_n268), .A3(new_n283), .A4(new_n266), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n266), .A2(new_n283), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n263), .A2(new_n269), .A3(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n282), .A2(new_n238), .A3(new_n284), .A4(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G902), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n188), .B1(new_n273), .B2(new_n289), .ZN(new_n290));
  AND2_X1   g104(.A1(new_n287), .A2(new_n288), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n239), .A2(new_n270), .A3(new_n272), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n291), .A2(new_n187), .A3(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G214), .B1(G237), .B2(G902), .ZN(new_n295));
  AOI21_X1  g109(.A(KEYINPUT80), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT80), .ZN(new_n297));
  INV_X1    g111(.A(new_n295), .ZN(new_n298));
  AOI211_X1 g112(.A(new_n297), .B(new_n298), .C1(new_n290), .C2(new_n293), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n205), .A2(G122), .ZN(new_n301));
  OR2_X1    g115(.A1(new_n301), .A2(KEYINPUT14), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(KEYINPUT14), .ZN(new_n303));
  INV_X1    g117(.A(G122), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G116), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G107), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n305), .A2(new_n301), .A3(new_n192), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n244), .A2(G128), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n250), .A2(G143), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G134), .B1(new_n311), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G134), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n310), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n307), .A2(new_n309), .A3(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT88), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT13), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT88), .A2(KEYINPUT13), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n313), .B1(new_n323), .B2(new_n311), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT89), .ZN(new_n325));
  AND2_X1   g139(.A1(KEYINPUT88), .A2(KEYINPUT13), .ZN(new_n326));
  NOR2_X1   g140(.A1(KEYINPUT88), .A2(KEYINPUT13), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n325), .B1(new_n328), .B2(new_n310), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n321), .A2(new_n310), .A3(new_n325), .A4(new_n322), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n324), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G134), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n192), .B1(new_n305), .B2(new_n301), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n316), .B1(new_n308), .B2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT90), .B1(new_n333), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT90), .ZN(new_n338));
  AOI211_X1 g152(.A(new_n338), .B(new_n335), .C1(new_n332), .C2(G134), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n318), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT9), .B(G234), .ZN(new_n341));
  INV_X1    g155(.A(G217), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n341), .A2(new_n342), .A3(G953), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT91), .ZN(new_n346));
  INV_X1    g160(.A(new_n318), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n321), .A2(new_n310), .A3(new_n322), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT89), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n330), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n315), .B1(new_n350), .B2(new_n324), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n338), .B1(new_n351), .B2(new_n335), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n312), .B1(new_n328), .B2(new_n310), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(new_n330), .B2(new_n349), .ZN(new_n354));
  OAI211_X1 g168(.A(KEYINPUT90), .B(new_n336), .C1(new_n354), .C2(new_n315), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n347), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n343), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n345), .A2(new_n346), .A3(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(KEYINPUT91), .A3(new_n343), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT92), .ZN(new_n361));
  INV_X1    g175(.A(G478), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(KEYINPUT15), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n360), .A2(new_n361), .A3(new_n288), .A4(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT20), .ZN(new_n366));
  NOR2_X1   g180(.A1(G475), .A2(G902), .ZN(new_n367));
  INV_X1    g181(.A(G237), .ZN(new_n368));
  INV_X1    g182(.A(G953), .ZN(new_n369));
  AND4_X1   g183(.A1(G143), .A2(new_n368), .A3(new_n369), .A4(G214), .ZN(new_n370));
  NOR2_X1   g184(.A1(G237), .A2(G953), .ZN(new_n371));
  AOI21_X1  g185(.A(G143), .B1(new_n371), .B2(G214), .ZN(new_n372));
  OAI21_X1  g186(.A(G131), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT17), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n368), .A2(new_n369), .A3(G214), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n244), .ZN(new_n376));
  INV_X1    g190(.A(G131), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n371), .A2(G143), .A3(G214), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n373), .A2(new_n374), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G125), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n254), .A2(G140), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(new_n383), .A3(KEYINPUT16), .ZN(new_n384));
  OR3_X1    g198(.A1(new_n254), .A2(KEYINPUT16), .A3(G140), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n242), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n384), .A2(new_n385), .A3(G146), .ZN(new_n388));
  OAI211_X1 g202(.A(KEYINPUT17), .B(G131), .C1(new_n370), .C2(new_n372), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n380), .A2(new_n387), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n382), .A2(new_n383), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G146), .ZN(new_n392));
  XNOR2_X1  g206(.A(G125), .B(G140), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n242), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n392), .A2(new_n394), .A3(KEYINPUT83), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT83), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n382), .A2(new_n383), .A3(new_n242), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n242), .B1(new_n382), .B2(new_n383), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(KEYINPUT82), .A2(KEYINPUT18), .A3(G131), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n370), .A2(new_n372), .A3(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n401), .B1(new_n376), .B2(new_n378), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g220(.A(G113), .B(G122), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT84), .B(G104), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n407), .A2(new_n408), .ZN(new_n411));
  OAI21_X1  g225(.A(KEYINPUT85), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n407), .A2(new_n408), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT85), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n414), .A3(new_n409), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n390), .A2(new_n406), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n413), .A2(new_n409), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n393), .A2(KEYINPUT19), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n393), .A2(KEYINPUT19), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n242), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n373), .A2(new_n379), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n388), .A2(KEYINPUT72), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT72), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n384), .A2(new_n385), .A3(new_n425), .A4(G146), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n422), .A2(new_n423), .A3(new_n424), .A4(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n418), .B1(new_n427), .B2(new_n406), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n366), .B(new_n367), .C1(new_n417), .C2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT86), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n390), .A2(new_n406), .A3(new_n416), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n393), .B(KEYINPUT19), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n432), .A2(new_n242), .B1(new_n373), .B2(new_n379), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n424), .A2(new_n426), .ZN(new_n434));
  AOI22_X1  g248(.A1(new_n433), .A2(new_n434), .B1(new_n400), .B2(new_n405), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n431), .B1(new_n435), .B2(new_n418), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n436), .A2(new_n437), .A3(new_n366), .A4(new_n367), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n367), .B1(new_n417), .B2(new_n428), .ZN(new_n439));
  XOR2_X1   g253(.A(KEYINPUT81), .B(KEYINPUT20), .Z(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n430), .A2(new_n438), .A3(new_n442), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n444), .A2(new_n380), .B1(new_n400), .B2(new_n405), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT87), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n418), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n390), .A2(new_n406), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT87), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n417), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G475), .B1(new_n450), .B2(G902), .ZN(new_n451));
  AND2_X1   g265(.A1(new_n369), .A2(G952), .ZN(new_n452));
  NAND2_X1  g266(.A1(G234), .A2(G237), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n454), .B(KEYINPUT93), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT21), .B(G898), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n453), .A2(G902), .A3(G953), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  AND3_X1   g273(.A1(new_n443), .A2(new_n451), .A3(new_n459), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n358), .A2(new_n361), .A3(new_n288), .A4(new_n359), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n363), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n365), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G469), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n315), .A2(G137), .ZN(new_n465));
  INV_X1    g279(.A(G137), .ZN(new_n466));
  AOI21_X1  g280(.A(KEYINPUT64), .B1(new_n466), .B2(G134), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT11), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n465), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT64), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n470), .B(new_n468), .C1(new_n315), .C2(G137), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(G131), .B1(new_n469), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n470), .B1(new_n315), .B2(G137), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT11), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n475), .A2(new_n377), .A3(new_n471), .A4(new_n465), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT12), .B1(new_n477), .B2(KEYINPUT78), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n201), .A2(new_n203), .ZN(new_n480));
  INV_X1    g294(.A(new_n267), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT75), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n246), .B2(new_n248), .ZN(new_n483));
  OAI211_X1 g297(.A(KEYINPUT75), .B(new_n247), .C1(new_n260), .C2(G128), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n252), .A3(new_n484), .ZN(new_n485));
  AOI22_X1  g299(.A1(new_n480), .A2(new_n481), .B1(new_n274), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n477), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n479), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n274), .ZN(new_n489));
  XNOR2_X1  g303(.A(KEYINPUT76), .B(KEYINPUT10), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n222), .A2(G101), .A3(new_n224), .ZN(new_n492));
  INV_X1    g306(.A(new_n231), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n264), .A3(new_n225), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n196), .A2(new_n199), .A3(new_n202), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n202), .B1(new_n196), .B2(new_n199), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n267), .A2(KEYINPUT10), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n491), .A2(new_n495), .A3(new_n487), .A4(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n489), .B1(new_n498), .B2(new_n267), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n477), .A3(new_n478), .ZN(new_n503));
  XNOR2_X1  g317(.A(G110), .B(G140), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n369), .A2(G227), .ZN(new_n505));
  XOR2_X1   g319(.A(new_n504), .B(new_n505), .Z(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n488), .A2(new_n501), .A3(new_n503), .A4(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n491), .A2(new_n495), .A3(new_n500), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n477), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n507), .B1(new_n511), .B2(new_n501), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n464), .B(new_n288), .C1(new_n509), .C2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n464), .A2(new_n288), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n488), .A2(new_n501), .A3(new_n503), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(new_n506), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n511), .A2(new_n501), .A3(new_n507), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(G469), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n513), .A2(new_n515), .A3(new_n519), .ZN(new_n520));
  OAI21_X1  g334(.A(G221), .B1(new_n341), .B2(G902), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g336(.A1(new_n463), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT32), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n371), .A2(G210), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT27), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT26), .B(G101), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT66), .ZN(new_n529));
  XNOR2_X1  g343(.A(new_n528), .B(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT65), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n229), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT65), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n476), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n466), .A2(G134), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n474), .B2(KEYINPUT11), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n377), .B1(new_n537), .B2(new_n471), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n264), .B1(new_n535), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n315), .A2(G137), .ZN(new_n540));
  OAI21_X1  g354(.A(G131), .B1(new_n540), .B2(new_n536), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n267), .A2(new_n476), .A3(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n534), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT28), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n539), .A2(new_n542), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n543), .A2(new_n544), .B1(new_n545), .B2(new_n229), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n534), .A2(new_n539), .A3(KEYINPUT28), .A4(new_n542), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n530), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n473), .A2(new_n476), .B1(new_n259), .B2(new_n261), .ZN(new_n549));
  AND3_X1   g363(.A1(new_n267), .A2(new_n476), .A3(new_n541), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT30), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT30), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n552), .B1(new_n539), .B2(new_n542), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n229), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(new_n543), .A3(new_n528), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT31), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n543), .ZN(new_n558));
  OAI21_X1  g372(.A(KEYINPUT30), .B1(new_n549), .B2(new_n550), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n539), .A2(new_n552), .A3(new_n542), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n558), .B1(new_n561), .B2(new_n229), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(KEYINPUT31), .A3(new_n528), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n548), .B1(new_n557), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(G472), .A2(G902), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT67), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n524), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n546), .A2(new_n547), .ZN(new_n568));
  INV_X1    g382(.A(new_n530), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT31), .B1(new_n562), .B2(new_n528), .ZN(new_n571));
  AOI22_X1  g385(.A1(new_n559), .A2(new_n560), .B1(new_n227), .B2(new_n228), .ZN(new_n572));
  INV_X1    g386(.A(new_n528), .ZN(new_n573));
  NOR4_X1   g387(.A1(new_n572), .A2(new_n558), .A3(new_n556), .A4(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n570), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n566), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(KEYINPUT32), .A3(new_n576), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n227), .A2(new_n228), .A3(KEYINPUT65), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT65), .B1(new_n227), .B2(new_n228), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n549), .B2(new_n550), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n581), .A2(new_n543), .A3(KEYINPUT68), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT68), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n545), .A2(new_n583), .A3(new_n580), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(KEYINPUT28), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n543), .A2(new_n544), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT29), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n573), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT69), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n589), .A2(new_n590), .A3(new_n288), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n589), .B2(new_n288), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n587), .B1(new_n562), .B2(new_n528), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n568), .A2(new_n569), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G472), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n567), .B(new_n577), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  OAI21_X1  g412(.A(KEYINPUT70), .B1(new_n250), .B2(G119), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT70), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n600), .A2(new_n209), .A3(G128), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n250), .A2(G119), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT24), .B(G110), .Z(new_n604));
  NAND2_X1  g418(.A1(new_n209), .A2(G128), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n250), .A2(KEYINPUT23), .A3(G119), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n209), .A2(G128), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(KEYINPUT23), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT71), .B(G110), .Z(new_n609));
  OAI22_X1  g423(.A1(new_n603), .A2(new_n604), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n610), .A2(new_n424), .A3(new_n426), .A4(new_n394), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n603), .A2(new_n604), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(G110), .ZN(new_n613));
  INV_X1    g427(.A(new_n388), .ZN(new_n614));
  AOI21_X1  g428(.A(G146), .B1(new_n384), .B2(new_n385), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n612), .B(new_n613), .C1(new_n614), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n611), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT22), .B(G137), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n369), .A2(G221), .A3(G234), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n611), .A2(new_n616), .A3(new_n620), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n288), .A3(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT25), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n622), .A2(KEYINPUT25), .A3(new_n288), .A4(new_n623), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n342), .B1(G234), .B2(new_n288), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT73), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n628), .A2(KEYINPUT73), .A3(new_n629), .ZN(new_n633));
  INV_X1    g447(.A(new_n623), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n620), .B1(new_n611), .B2(new_n616), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n629), .A2(G902), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n632), .A2(new_n633), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n300), .A2(new_n523), .A3(new_n598), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G101), .ZN(G3));
  INV_X1    g456(.A(KEYINPUT94), .ZN(new_n643));
  OAI21_X1  g457(.A(G472), .B1(new_n564), .B2(G902), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT73), .B1(new_n628), .B2(new_n629), .ZN(new_n645));
  INV_X1    g459(.A(new_n629), .ZN(new_n646));
  AOI211_X1 g460(.A(new_n631), .B(new_n646), .C1(new_n626), .C2(new_n627), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n575), .A2(new_n576), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n644), .A2(new_n648), .A3(new_n649), .A4(new_n638), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n643), .B1(new_n650), .B2(new_n522), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n597), .B1(new_n575), .B2(new_n288), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n564), .A2(new_n566), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n521), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n489), .A2(new_n490), .B1(new_n498), .B2(new_n499), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n487), .B1(new_n656), .B2(new_n495), .ZN(new_n657));
  AND4_X1   g471(.A1(new_n487), .A2(new_n491), .A3(new_n495), .A4(new_n500), .ZN(new_n658));
  OAI21_X1  g472(.A(new_n506), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(G902), .B1(new_n659), .B2(new_n508), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n514), .B1(new_n660), .B2(new_n464), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n655), .B1(new_n661), .B2(new_n519), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n654), .A2(new_n662), .A3(new_n640), .A4(KEYINPUT94), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n651), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n443), .A2(new_n451), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT95), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n340), .A2(new_n667), .A3(new_n344), .ZN(new_n668));
  OAI21_X1  g482(.A(KEYINPUT95), .B1(new_n356), .B2(new_n343), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT33), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n356), .B2(new_n343), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n668), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(KEYINPUT96), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT96), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n668), .A2(new_n669), .A3(new_n671), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n358), .A2(new_n670), .A3(new_n359), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n362), .A2(G902), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n676), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n358), .A2(new_n288), .A3(new_n359), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n362), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n666), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  AOI211_X1 g496(.A(new_n298), .B(new_n458), .C1(new_n290), .C2(new_n293), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n664), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT34), .B(G104), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G6));
  INV_X1    g501(.A(new_n451), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n439), .A2(new_n441), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n440), .B1(new_n436), .B2(new_n367), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT97), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n690), .A2(new_n691), .A3(KEYINPUT98), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT98), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n442), .B2(KEYINPUT97), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n689), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(KEYINPUT98), .B1(new_n690), .B2(new_n691), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n442), .A2(KEYINPUT97), .A3(new_n693), .ZN(new_n697));
  INV_X1    g511(.A(new_n689), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n688), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n365), .A2(new_n462), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n683), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n664), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT35), .B(G107), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G9));
  NOR2_X1   g519(.A1(new_n621), .A2(KEYINPUT36), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n617), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n637), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n632), .A2(new_n633), .A3(new_n708), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n709), .A2(new_n644), .A3(new_n649), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n300), .A2(new_n523), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT37), .B(G110), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G12));
  AND3_X1   g527(.A1(new_n632), .A2(new_n633), .A3(new_n708), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n273), .A2(new_n188), .A3(new_n289), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n187), .B1(new_n291), .B2(new_n292), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n295), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n522), .A2(new_n714), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(G900), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n455), .B1(new_n719), .B2(new_n457), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n698), .B1(new_n696), .B2(new_n697), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n451), .B(new_n721), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n461), .B(new_n364), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n718), .A2(new_n598), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G128), .ZN(G30));
  XOR2_X1   g542(.A(new_n720), .B(KEYINPUT39), .Z(new_n729));
  NAND2_X1  g543(.A1(new_n662), .A2(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(new_n730), .B(KEYINPUT40), .Z(new_n731));
  XOR2_X1   g545(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n732));
  XNOR2_X1  g546(.A(new_n294), .B(new_n732), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n733), .A2(new_n298), .A3(new_n709), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n701), .A2(new_n665), .ZN(new_n735));
  NOR3_X1   g549(.A1(new_n564), .A2(new_n524), .A3(new_n566), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT32), .B1(new_n575), .B2(new_n576), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT100), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n569), .A2(new_n584), .A3(new_n582), .ZN(new_n740));
  INV_X1    g554(.A(new_n555), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n288), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(G472), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n738), .A2(new_n739), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n567), .A2(new_n577), .A3(new_n743), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT100), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n735), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n731), .A2(new_n734), .A3(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G143), .ZN(G45));
  AOI211_X1 g563(.A(new_n666), .B(new_n720), .C1(new_n679), .C2(new_n681), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n718), .A2(new_n750), .A3(new_n598), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G146), .ZN(G48));
  OAI21_X1  g566(.A(new_n288), .B1(new_n509), .B2(new_n512), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(G469), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n521), .A3(new_n513), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n592), .A2(new_n595), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n589), .A2(new_n590), .A3(new_n288), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n597), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n567), .A2(new_n577), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n756), .B(new_n640), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n684), .ZN(new_n762));
  XOR2_X1   g576(.A(KEYINPUT41), .B(G113), .Z(new_n763));
  XNOR2_X1  g577(.A(new_n762), .B(new_n763), .ZN(G15));
  NOR2_X1   g578(.A1(new_n761), .A2(new_n702), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n205), .ZN(G18));
  INV_X1    g580(.A(KEYINPUT101), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n767), .B1(new_n755), .B2(new_n717), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n659), .A2(new_n508), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n464), .B1(new_n769), .B2(new_n288), .ZN(new_n770));
  AOI211_X1 g584(.A(G469), .B(G902), .C1(new_n659), .C2(new_n508), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n298), .B1(new_n290), .B2(new_n293), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n772), .A2(KEYINPUT101), .A3(new_n773), .A4(new_n521), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n589), .A2(new_n288), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(KEYINPUT69), .ZN(new_n777));
  OR2_X1    g591(.A1(new_n593), .A2(new_n594), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n777), .A2(new_n778), .A3(new_n758), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(G472), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n714), .B1(new_n738), .B2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n463), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n775), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT102), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n775), .A2(new_n781), .A3(KEYINPUT102), .A4(new_n782), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G119), .ZN(G21));
  NOR2_X1   g602(.A1(new_n725), .A2(new_n666), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n557), .A2(new_n563), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n585), .A2(new_n586), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n569), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n566), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n639), .A2(new_n652), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n755), .A2(new_n458), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n789), .A2(new_n794), .A3(new_n773), .A4(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G122), .ZN(G24));
  NOR3_X1   g611(.A1(new_n714), .A2(new_n652), .A3(new_n793), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n775), .A2(new_n750), .A3(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G125), .ZN(G27));
  NAND3_X1  g614(.A1(new_n682), .A2(KEYINPUT42), .A3(new_n721), .ZN(new_n801));
  AND3_X1   g615(.A1(new_n516), .A2(KEYINPUT103), .A3(new_n506), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT103), .B1(new_n516), .B2(new_n506), .ZN(new_n803));
  OAI211_X1 g617(.A(G469), .B(new_n518), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n655), .B1(new_n661), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT104), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n290), .A2(new_n295), .A3(new_n293), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n810), .B1(new_n805), .B2(new_n806), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n801), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  AOI22_X1  g626(.A1(G472), .A2(new_n779), .B1(new_n567), .B2(KEYINPUT105), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT105), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n814), .B1(new_n736), .B2(new_n737), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n639), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n816), .A2(KEYINPUT106), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT106), .ZN(new_n818));
  AOI211_X1 g632(.A(new_n818), .B(new_n639), .C1(new_n813), .C2(new_n815), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n812), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n661), .A2(new_n804), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n521), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n809), .B1(new_n822), .B2(KEYINPUT104), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n639), .B1(new_n738), .B2(new_n780), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n824), .A3(new_n750), .A4(new_n807), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT42), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n820), .A2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(G131), .ZN(G33));
  NAND4_X1  g643(.A1(new_n823), .A2(new_n824), .A3(new_n726), .A4(new_n807), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G134), .ZN(G36));
  AOI22_X1  g645(.A1(new_n670), .A2(new_n360), .B1(new_n673), .B2(new_n675), .ZN(new_n832));
  AOI22_X1  g646(.A1(new_n832), .A2(new_n678), .B1(new_n362), .B2(new_n680), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(new_n665), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT43), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n654), .A2(new_n714), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n835), .A2(KEYINPUT44), .A3(new_n836), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n837), .A2(new_n810), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT45), .B1(new_n517), .B2(new_n518), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n464), .ZN(new_n840));
  OAI211_X1 g654(.A(KEYINPUT45), .B(new_n518), .C1(new_n802), .C2(new_n803), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(new_n515), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT46), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n771), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(new_n844), .B2(new_n843), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n521), .A3(new_n729), .ZN(new_n847));
  OR2_X1    g661(.A1(new_n847), .A2(KEYINPUT107), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(KEYINPUT107), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n835), .A2(new_n836), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT44), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n838), .A2(new_n850), .A3(new_n853), .ZN(new_n854));
  XOR2_X1   g668(.A(KEYINPUT108), .B(G137), .Z(new_n855));
  XNOR2_X1  g669(.A(new_n854), .B(new_n855), .ZN(G39));
  NOR3_X1   g670(.A1(new_n598), .A2(new_n640), .A3(new_n809), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n846), .A2(KEYINPUT47), .A3(new_n521), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  AOI21_X1  g673(.A(KEYINPUT47), .B1(new_n846), .B2(new_n521), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n750), .B(new_n857), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(G140), .ZN(G42));
  NAND4_X1  g676(.A1(new_n823), .A2(new_n750), .A3(new_n798), .A4(new_n807), .ZN(new_n863));
  OAI21_X1  g677(.A(KEYINPUT111), .B1(new_n724), .B2(new_n701), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT111), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n700), .A2(new_n725), .A3(new_n865), .A4(new_n721), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n522), .A2(new_n809), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n781), .A2(new_n864), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n830), .A2(new_n863), .A3(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n823), .A2(KEYINPUT42), .A3(new_n750), .A4(new_n807), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n596), .A2(new_n597), .B1(new_n737), .B2(new_n814), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT105), .B1(new_n567), .B2(new_n577), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n640), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(new_n818), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n816), .A2(KEYINPUT106), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n870), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n825), .A2(new_n826), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n869), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n641), .A2(new_n711), .A3(new_n796), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n761), .B1(new_n684), .B2(new_n702), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT109), .B1(new_n833), .B2(new_n666), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT109), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n682), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT110), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n886), .B1(new_n725), .B2(new_n665), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n701), .A2(KEYINPUT110), .A3(new_n666), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n296), .A2(new_n299), .A3(new_n458), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(new_n651), .A3(new_n663), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n890), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n881), .A2(new_n787), .A3(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n878), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT52), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n598), .B(new_n718), .C1(new_n750), .C2(new_n726), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n799), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n745), .B(new_n739), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n900), .A2(new_n717), .A3(new_n735), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n720), .B(KEYINPUT112), .Z(new_n902));
  NAND4_X1  g716(.A1(new_n632), .A2(new_n633), .A3(new_n708), .A4(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT113), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT113), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n648), .A2(new_n905), .A3(new_n708), .A4(new_n902), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT114), .B1(new_n907), .B2(new_n805), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n907), .A2(KEYINPUT114), .A3(new_n805), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n899), .B1(new_n901), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n897), .B1(new_n912), .B2(KEYINPUT115), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n898), .A2(new_n799), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n907), .A2(KEYINPUT114), .A3(new_n805), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n773), .B(new_n747), .C1(new_n915), .C2(new_n908), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT115), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n918), .A3(KEYINPUT52), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n896), .A2(new_n913), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT53), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n920), .A2(KEYINPUT116), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(KEYINPUT52), .B1(new_n914), .B2(new_n916), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n914), .A2(new_n916), .A3(KEYINPUT52), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n896), .B(KEYINPUT53), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT116), .B1(new_n920), .B2(new_n921), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT54), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n924), .A2(new_n923), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n830), .A2(new_n863), .A3(new_n868), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n930), .B1(new_n820), .B2(new_n827), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n679), .A2(new_n681), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n932), .A2(new_n665), .A3(new_n683), .ZN(new_n933));
  AND3_X1   g747(.A1(new_n683), .A2(new_n700), .A3(new_n701), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n824), .B(new_n756), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n935), .A2(new_n641), .A3(new_n711), .A4(new_n796), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n892), .B1(new_n885), .B2(new_n889), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g752(.A1(new_n931), .A2(new_n938), .A3(new_n787), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n921), .B1(new_n929), .B2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n896), .A2(KEYINPUT53), .A3(new_n913), .A4(new_n919), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT54), .ZN(new_n942));
  AND3_X1   g756(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n928), .A2(new_n944), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n835), .A2(new_n455), .A3(new_n794), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT50), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n295), .B1(KEYINPUT118), .B2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n733), .A2(new_n756), .A3(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n947), .A2(KEYINPUT118), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n835), .A2(new_n455), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n755), .A2(new_n809), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n798), .A3(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n900), .A2(new_n640), .A3(new_n455), .A4(new_n955), .ZN(new_n957));
  OR3_X1    g771(.A1(new_n957), .A2(new_n665), .A3(new_n932), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n953), .A2(new_n956), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n859), .A2(new_n860), .ZN(new_n960));
  OR2_X1    g774(.A1(new_n772), .A2(KEYINPUT117), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n772), .A2(KEYINPUT117), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n961), .A2(new_n655), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  AND3_X1   g778(.A1(new_n964), .A2(new_n810), .A3(new_n946), .ZN(new_n965));
  INV_X1    g779(.A(new_n965), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n951), .A2(new_n952), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n959), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT51), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n959), .A2(new_n966), .A3(KEYINPUT51), .A4(new_n967), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n946), .A2(new_n775), .ZN(new_n972));
  INV_X1    g786(.A(new_n682), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n972), .B(new_n452), .C1(new_n973), .C2(new_n957), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n874), .A2(new_n875), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n954), .A2(new_n975), .A3(new_n955), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(KEYINPUT48), .ZN(new_n977));
  OR2_X1    g791(.A1(new_n976), .A2(KEYINPUT48), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n970), .A2(new_n971), .A3(new_n979), .ZN(new_n980));
  OAI22_X1  g794(.A1(new_n945), .A2(new_n980), .B1(G952), .B2(G953), .ZN(new_n981));
  AND4_X1   g795(.A1(new_n640), .A2(new_n733), .A3(new_n295), .A4(new_n521), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n772), .B(KEYINPUT49), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n982), .A2(new_n900), .A3(new_n834), .A4(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n981), .A2(new_n984), .ZN(G75));
  NOR2_X1   g799(.A1(new_n369), .A2(G952), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n288), .B1(new_n940), .B2(new_n941), .ZN(new_n988));
  AOI21_X1  g802(.A(KEYINPUT56), .B1(new_n988), .B2(G210), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n239), .A2(new_n272), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(new_n270), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT55), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n987), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n989), .B2(new_n993), .ZN(G51));
  AOI211_X1 g809(.A(new_n288), .B(new_n842), .C1(new_n940), .C2(new_n941), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n514), .B(KEYINPUT57), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n942), .B1(new_n940), .B2(new_n941), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n997), .B1(new_n943), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n769), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT119), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n996), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n999), .A2(KEYINPUT119), .A3(new_n769), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n986), .B1(new_n1002), .B2(new_n1003), .ZN(G54));
  NAND3_X1  g818(.A1(new_n988), .A2(KEYINPUT58), .A3(G475), .ZN(new_n1005));
  INV_X1    g819(.A(new_n436), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n1005), .A2(KEYINPUT120), .A3(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n987), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1008));
  AOI21_X1  g822(.A(KEYINPUT120), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(G60));
  XOR2_X1   g824(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1011));
  NOR2_X1   g825(.A1(new_n362), .A2(new_n288), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1011), .B(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n832), .B1(new_n945), .B2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n832), .B(new_n1014), .C1(new_n943), .C2(new_n998), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1016), .A2(new_n987), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n1015), .A2(new_n1017), .ZN(G63));
  NAND2_X1  g832(.A1(new_n940), .A2(new_n941), .ZN(new_n1019));
  XNOR2_X1  g833(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n342), .A2(new_n288), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1019), .A2(new_n707), .A3(new_n1022), .ZN(new_n1023));
  NOR2_X1   g837(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n986), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n636), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g842(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n1029));
  XOR2_X1   g843(.A(new_n1029), .B(KEYINPUT124), .Z(new_n1030));
  XNOR2_X1  g844(.A(new_n1028), .B(new_n1030), .ZN(G66));
  NOR3_X1   g845(.A1(new_n456), .A2(new_n240), .A3(new_n369), .ZN(new_n1032));
  INV_X1    g846(.A(new_n895), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1032), .B1(new_n1033), .B2(new_n369), .ZN(new_n1034));
  INV_X1    g848(.A(G898), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n990), .B1(new_n1035), .B2(G953), .ZN(new_n1036));
  XOR2_X1   g850(.A(new_n1034), .B(new_n1036), .Z(G69));
  NAND2_X1  g851(.A1(new_n748), .A2(new_n914), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT62), .ZN(new_n1039));
  XNOR2_X1  g853(.A(new_n1038), .B(new_n1039), .ZN(new_n1040));
  NOR2_X1   g854(.A1(new_n730), .A2(new_n809), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n890), .A2(new_n824), .A3(new_n1041), .ZN(new_n1042));
  NAND4_X1  g856(.A1(new_n1040), .A2(new_n854), .A3(new_n861), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(new_n369), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n561), .B(new_n432), .Z(new_n1045));
  NAND2_X1  g859(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1045), .B1(G900), .B2(G953), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n853), .A2(new_n810), .A3(new_n837), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n735), .A2(new_n717), .ZN(new_n1049));
  NAND2_X1  g863(.A1(new_n975), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1051), .A2(new_n850), .ZN(new_n1052));
  AND3_X1   g866(.A1(new_n828), .A2(new_n830), .A3(new_n914), .ZN(new_n1053));
  AND2_X1   g867(.A1(new_n1053), .A2(new_n861), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g869(.A(new_n1047), .B1(new_n1055), .B2(G953), .ZN(new_n1056));
  INV_X1    g870(.A(KEYINPUT125), .ZN(new_n1057));
  NAND3_X1  g871(.A1(new_n1046), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1047), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1053), .A2(new_n861), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n1060), .B1(new_n850), .B2(new_n1051), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n1059), .B1(new_n1061), .B2(new_n369), .ZN(new_n1062));
  INV_X1    g876(.A(new_n1045), .ZN(new_n1063));
  AOI21_X1  g877(.A(new_n1063), .B1(new_n1043), .B2(new_n369), .ZN(new_n1064));
  OAI21_X1  g878(.A(KEYINPUT125), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g879(.A(new_n369), .B1(G227), .B2(G900), .ZN(new_n1066));
  AND3_X1   g880(.A1(new_n1058), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  AOI21_X1  g881(.A(new_n1066), .B1(new_n1058), .B2(new_n1065), .ZN(new_n1068));
  NOR2_X1   g882(.A1(new_n1067), .A2(new_n1068), .ZN(G72));
  NAND2_X1  g883(.A1(G472), .A2(G902), .ZN(new_n1070));
  XOR2_X1   g884(.A(new_n1070), .B(KEYINPUT63), .Z(new_n1071));
  OAI21_X1  g885(.A(new_n1071), .B1(new_n1055), .B2(new_n895), .ZN(new_n1072));
  NOR3_X1   g886(.A1(new_n572), .A2(new_n558), .A3(new_n528), .ZN(new_n1073));
  NAND2_X1  g887(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  OAI21_X1  g888(.A(new_n1071), .B1(new_n1043), .B2(new_n895), .ZN(new_n1075));
  NOR2_X1   g889(.A1(new_n562), .A2(new_n573), .ZN(new_n1076));
  NAND2_X1  g890(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g891(.A1(new_n1074), .A2(new_n1077), .A3(new_n987), .ZN(new_n1078));
  INV_X1    g892(.A(new_n1071), .ZN(new_n1079));
  NOR3_X1   g893(.A1(new_n1076), .A2(new_n1073), .A3(new_n1079), .ZN(new_n1080));
  XOR2_X1   g894(.A(new_n1080), .B(KEYINPUT126), .Z(new_n1081));
  OAI21_X1  g895(.A(new_n1081), .B1(new_n926), .B2(new_n927), .ZN(new_n1082));
  OR2_X1    g896(.A1(new_n1082), .A2(KEYINPUT127), .ZN(new_n1083));
  NAND2_X1  g897(.A1(new_n1082), .A2(KEYINPUT127), .ZN(new_n1084));
  AOI21_X1  g898(.A(new_n1078), .B1(new_n1083), .B2(new_n1084), .ZN(G57));
endmodule


