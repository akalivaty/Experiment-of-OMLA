//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 0 1 0 0 0 0 0 1 1 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n697, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G953), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT70), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT70), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G953), .ZN(new_n196));
  AND2_X1   g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G227), .ZN(new_n198));
  XOR2_X1   g012(.A(G110), .B(G140), .Z(new_n199));
  XNOR2_X1  g013(.A(new_n198), .B(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI211_X1 g019(.A(KEYINPUT67), .B(KEYINPUT1), .C1(new_n203), .C2(G146), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G128), .ZN(new_n207));
  AOI21_X1  g021(.A(KEYINPUT67), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n205), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT65), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n210), .B1(new_n203), .B2(G146), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n201), .A2(KEYINPUT65), .A3(G143), .ZN(new_n212));
  INV_X1    g026(.A(G128), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(KEYINPUT1), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n211), .A2(new_n212), .A3(new_n214), .A4(new_n204), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n209), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G104), .ZN(new_n217));
  NOR3_X1   g031(.A1(new_n217), .A2(KEYINPUT3), .A3(G107), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT75), .B(G104), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n218), .B1(new_n219), .B2(G107), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n217), .A2(KEYINPUT75), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT75), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G104), .ZN(new_n225));
  AOI21_X1  g039(.A(G107), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n220), .B(new_n221), .C1(new_n222), .C2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G107), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(G104), .ZN(new_n229));
  OAI21_X1  g043(.A(G101), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n216), .A2(new_n227), .A3(KEYINPUT10), .A4(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n231), .B(KEYINPUT76), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT11), .ZN(new_n233));
  INV_X1    g047(.A(G134), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(G137), .ZN(new_n235));
  INV_X1    g049(.A(G137), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT11), .A3(G134), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(G137), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G131), .ZN(new_n240));
  INV_X1    g054(.A(G131), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n235), .A2(new_n237), .A3(new_n241), .A4(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n223), .A2(new_n225), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n222), .B1(new_n244), .B2(new_n228), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n223), .A2(new_n225), .A3(G107), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n222), .A2(new_n228), .A3(G104), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g062(.A(G101), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n227), .A2(new_n249), .A3(KEYINPUT4), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n211), .A2(new_n212), .A3(new_n204), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(KEYINPUT0), .A2(G128), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n254), .B1(new_n202), .B2(new_n204), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT0), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(new_n213), .A3(KEYINPUT64), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT64), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(KEYINPUT0), .B2(G128), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n252), .A2(new_n254), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n262), .B(G101), .C1(new_n245), .C2(new_n248), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n250), .A2(new_n261), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n213), .B1(new_n202), .B2(KEYINPUT1), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n215), .B1(new_n252), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n227), .A2(new_n266), .A3(new_n230), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT10), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n264), .A2(new_n269), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n232), .A2(new_n243), .A3(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(new_n240), .A2(new_n242), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n264), .A2(new_n269), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT76), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n231), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n244), .A2(new_n228), .ZN(new_n276));
  INV_X1    g090(.A(new_n229), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n221), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n245), .A2(new_n248), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n278), .B1(new_n279), .B2(new_n221), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n280), .A2(KEYINPUT76), .A3(KEYINPUT10), .A4(new_n216), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n272), .B1(new_n273), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n200), .B1(new_n271), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n267), .B1(new_n280), .B2(new_n216), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT12), .ZN(new_n286));
  AND2_X1   g100(.A1(new_n243), .A2(KEYINPUT77), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n286), .B1(new_n285), .B2(new_n287), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n282), .A2(new_n272), .A3(new_n269), .A4(new_n264), .ZN(new_n292));
  INV_X1    g106(.A(new_n200), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n284), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n192), .B1(new_n295), .B2(new_n190), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n292), .A2(new_n293), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n297), .A2(new_n283), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n293), .B1(new_n291), .B2(new_n292), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT78), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n290), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n288), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n200), .B1(new_n271), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT78), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n243), .B1(new_n232), .B2(new_n270), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n292), .A3(new_n293), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n300), .A2(new_n307), .A3(G469), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n189), .B1(new_n296), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(G214), .B1(G237), .B2(G902), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(KEYINPUT79), .ZN(new_n311));
  OAI21_X1  g125(.A(G210), .B1(G237), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G116), .ZN(new_n314));
  OAI21_X1  g128(.A(KEYINPUT68), .B1(new_n314), .B2(G119), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT68), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n316), .A2(new_n317), .A3(G116), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n314), .A2(G119), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n315), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G113), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(KEYINPUT2), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT2), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G113), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n315), .A2(new_n318), .A3(KEYINPUT5), .A4(new_n319), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n314), .A2(KEYINPUT5), .A3(G119), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(new_n322), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n321), .A2(new_n326), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n280), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n250), .A2(new_n263), .ZN(new_n332));
  INV_X1    g146(.A(new_n326), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n320), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n326), .A2(new_n315), .A3(new_n318), .A4(new_n319), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n334), .A2(KEYINPUT69), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT69), .B1(new_n334), .B2(new_n335), .ZN(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n331), .B1(new_n332), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(G110), .B(G122), .ZN(new_n340));
  XOR2_X1   g154(.A(new_n340), .B(KEYINPUT80), .Z(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n339), .A2(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n341), .B(new_n331), .C1(new_n332), .C2(new_n338), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(KEYINPUT6), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n260), .A2(new_n205), .A3(new_n253), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n251), .B2(new_n253), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(G125), .ZN(new_n348));
  INV_X1    g162(.A(G125), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n209), .A2(new_n349), .A3(new_n215), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n193), .A2(G224), .ZN(new_n352));
  XOR2_X1   g166(.A(new_n352), .B(KEYINPUT81), .Z(new_n353));
  XOR2_X1   g167(.A(new_n351), .B(new_n353), .Z(new_n354));
  INV_X1    g168(.A(KEYINPUT6), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n339), .A2(new_n355), .A3(new_n342), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n345), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(new_n191), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT82), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n227), .B(new_n230), .C1(new_n330), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n327), .A2(new_n329), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n335), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(KEYINPUT82), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT83), .B1(new_n360), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n330), .A2(new_n359), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n362), .A2(KEYINPUT82), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT83), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n280), .A2(new_n365), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  OR2_X1    g182(.A1(new_n280), .A2(new_n330), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n364), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n341), .B(KEYINPUT8), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n370), .A2(KEYINPUT84), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(KEYINPUT84), .B1(new_n370), .B2(new_n371), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n348), .A2(KEYINPUT7), .A3(new_n353), .A4(new_n350), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n348), .A2(new_n350), .B1(KEYINPUT7), .B2(new_n353), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n375), .A2(KEYINPUT85), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT85), .ZN(new_n377));
  AOI221_X4 g191(.A(new_n377), .B1(KEYINPUT7), .B2(new_n353), .C1(new_n348), .C2(new_n350), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n344), .B(new_n374), .C1(new_n376), .C2(new_n378), .ZN(new_n379));
  NOR3_X1   g193(.A1(new_n372), .A2(new_n373), .A3(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n313), .B1(new_n358), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n379), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n370), .A2(new_n371), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n370), .A2(KEYINPUT84), .A3(new_n371), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n387), .A2(new_n191), .A3(new_n312), .A4(new_n357), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n311), .B1(new_n381), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G217), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n187), .A2(new_n390), .A3(G953), .ZN(new_n391));
  INV_X1    g205(.A(G122), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G116), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n392), .A2(G116), .ZN(new_n395));
  OAI21_X1  g209(.A(G107), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n395), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n397), .A2(new_n228), .A3(new_n393), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n213), .A2(G143), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n203), .A2(G128), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n396), .A2(new_n398), .B1(new_n234), .B2(new_n401), .ZN(new_n402));
  XOR2_X1   g216(.A(KEYINPUT86), .B(KEYINPUT13), .Z(new_n403));
  INV_X1    g217(.A(new_n399), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT87), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n400), .B1(new_n403), .B2(new_n404), .ZN(new_n406));
  XNOR2_X1  g220(.A(KEYINPUT86), .B(KEYINPUT13), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(new_n399), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n405), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT88), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n410), .A2(new_n411), .A3(G134), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n411), .B1(new_n410), .B2(G134), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n402), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n401), .B(new_n234), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT89), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n416), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT14), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n395), .B1(new_n419), .B2(new_n393), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT90), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n228), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT90), .B1(new_n397), .B2(KEYINPUT14), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n422), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n417), .A2(new_n418), .A3(new_n398), .A4(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n391), .B1(new_n414), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n414), .A2(new_n425), .A3(new_n391), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n191), .ZN(new_n430));
  INV_X1    g244(.A(G478), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n431), .A2(KEYINPUT15), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n429), .B(new_n191), .C1(KEYINPUT15), .C2(new_n431), .ZN(new_n434));
  INV_X1    g248(.A(new_n197), .ZN(new_n435));
  NAND2_X1  g249(.A1(G234), .A2(G237), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n435), .A2(G902), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(G898), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n436), .A2(G952), .A3(new_n193), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n433), .A2(new_n434), .A3(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(G113), .B(G122), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(new_n217), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G237), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n194), .A2(new_n196), .A3(G214), .A4(new_n447), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n448), .A2(new_n203), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n203), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT18), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(new_n241), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(G125), .B(G140), .ZN(new_n455));
  XNOR2_X1  g269(.A(new_n455), .B(new_n201), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n449), .B(new_n450), .C1(new_n452), .C2(new_n241), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n455), .A2(KEYINPUT16), .ZN(new_n460));
  OR3_X1    g274(.A1(new_n349), .A2(KEYINPUT16), .A3(G140), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(G146), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT73), .ZN(new_n463));
  AND2_X1   g277(.A1(new_n455), .A2(KEYINPUT19), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n455), .A2(KEYINPUT19), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n201), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT73), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n460), .A2(new_n467), .A3(new_n461), .A4(G146), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n463), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n449), .A2(new_n241), .A3(new_n450), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n451), .A2(G131), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n446), .B1(new_n459), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT17), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n471), .A2(new_n474), .A3(new_n470), .ZN(new_n475));
  INV_X1    g289(.A(new_n462), .ZN(new_n476));
  AOI21_X1  g290(.A(G146), .B1(new_n460), .B2(new_n461), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(new_n471), .B2(new_n474), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n445), .B(new_n458), .C1(new_n475), .C2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n473), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT20), .ZN(new_n482));
  NOR2_X1   g296(.A1(G475), .A2(G902), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n482), .B1(new_n481), .B2(new_n483), .ZN(new_n486));
  INV_X1    g300(.A(G475), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n458), .B1(new_n475), .B2(new_n479), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n446), .ZN(new_n489));
  AOI21_X1  g303(.A(G902), .B1(new_n489), .B2(new_n480), .ZN(new_n490));
  OAI22_X1  g304(.A1(new_n485), .A2(new_n486), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n443), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n309), .A2(new_n389), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT91), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT32), .ZN(new_n496));
  INV_X1    g310(.A(new_n238), .ZN(new_n497));
  NOR2_X1   g311(.A1(new_n234), .A2(G137), .ZN(new_n498));
  OAI21_X1  g312(.A(G131), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n499), .A2(new_n242), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n216), .A2(new_n501), .B1(new_n261), .B2(new_n243), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT28), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n502), .A2(new_n338), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n503), .B1(new_n502), .B2(new_n338), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n500), .B1(new_n209), .B2(new_n215), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT66), .B1(new_n272), .B2(new_n347), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT66), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n261), .A2(new_n243), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n506), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n504), .A2(new_n505), .B1(new_n510), .B2(new_n338), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n197), .A2(G210), .A3(new_n447), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT27), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT26), .B(G101), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n338), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n502), .A2(KEYINPUT30), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n518), .B(new_n519), .C1(new_n510), .C2(KEYINPUT30), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT31), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n502), .A2(new_n338), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n520), .A2(new_n521), .A3(new_n515), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n520), .A2(new_n515), .A3(new_n522), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT31), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT71), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT71), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n528), .A3(KEYINPUT31), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n524), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(G472), .A2(G902), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n496), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n502), .A2(new_n338), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n535), .B1(new_n504), .B2(new_n505), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n515), .A2(KEYINPUT29), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n520), .A2(new_n522), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(new_n515), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT29), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n540), .B1(new_n511), .B2(new_n516), .ZN(new_n541));
  OAI221_X1 g355(.A(new_n191), .B1(new_n536), .B2(new_n537), .C1(new_n539), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G472), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n517), .A2(new_n523), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n525), .A2(new_n528), .A3(KEYINPUT31), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n528), .B1(new_n525), .B2(KEYINPUT31), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n547), .A2(KEYINPUT32), .A3(new_n531), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n533), .A2(new_n543), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n390), .B1(G234), .B2(new_n191), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n213), .A2(G119), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n317), .A2(G128), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  XNOR2_X1  g367(.A(KEYINPUT24), .B(G110), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT72), .ZN(new_n556));
  INV_X1    g370(.A(G110), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT23), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n213), .A2(KEYINPUT23), .A3(G119), .ZN(new_n560));
  AND3_X1   g374(.A1(new_n559), .A2(new_n560), .A3(new_n552), .ZN(new_n561));
  OAI221_X1 g375(.A(new_n556), .B1(new_n557), .B2(new_n561), .C1(new_n477), .C2(new_n476), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n561), .A2(new_n557), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n553), .A2(new_n554), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n563), .A2(new_n564), .B1(new_n201), .B2(new_n455), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(new_n463), .A3(new_n468), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT74), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n562), .A2(KEYINPUT74), .A3(new_n566), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n197), .A2(G221), .A3(G234), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT22), .B(G137), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n571), .B(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n569), .A2(new_n570), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n567), .A2(new_n568), .A3(new_n573), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND3_X1   g391(.A1(new_n577), .A2(KEYINPUT25), .A3(new_n191), .ZN(new_n578));
  AOI21_X1  g392(.A(KEYINPUT25), .B1(new_n577), .B2(new_n191), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n550), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n550), .A2(G902), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n549), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n309), .A2(KEYINPUT91), .A3(new_n389), .A4(new_n492), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n495), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n428), .B2(KEYINPUT94), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT94), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n414), .A2(new_n592), .A3(new_n425), .A4(new_n391), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT93), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n426), .A2(new_n594), .ZN(new_n595));
  AOI211_X1 g409(.A(KEYINPUT93), .B(new_n391), .C1(new_n414), .C2(new_n425), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n591), .B(new_n593), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n429), .A2(new_n590), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n431), .A2(G902), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(KEYINPUT95), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n430), .A2(new_n431), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT95), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n597), .A2(new_n598), .A3(new_n603), .A4(new_n599), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n601), .A2(new_n602), .A3(new_n604), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n605), .A2(new_n491), .A3(new_n442), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT92), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n388), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n381), .ZN(new_n609));
  OAI211_X1 g423(.A(new_n607), .B(new_n313), .C1(new_n358), .C2(new_n380), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n311), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n606), .A2(new_n611), .ZN(new_n612));
  OAI21_X1  g426(.A(G472), .B1(new_n530), .B2(G902), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n547), .A2(new_n531), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n616), .A2(new_n584), .A3(new_n309), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT34), .B(G104), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  INV_X1    g434(.A(new_n617), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n485), .A2(new_n486), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT96), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n490), .A2(new_n487), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n433), .A2(new_n434), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n442), .B(KEYINPUT97), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  AOI211_X1 g443(.A(new_n311), .B(new_n629), .C1(new_n609), .C2(new_n610), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n621), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n631), .B(KEYINPUT98), .Z(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NOR2_X1   g448(.A1(new_n574), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n567), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n581), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n580), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n615), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n495), .A2(new_n587), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT37), .B(G110), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(G12));
  INV_X1    g457(.A(G900), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n440), .B1(new_n437), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n627), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n611), .A2(new_n549), .A3(new_n309), .A4(new_n638), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n213), .ZN(G30));
  INV_X1    g464(.A(new_n533), .ZN(new_n651));
  INV_X1    g465(.A(new_n548), .ZN(new_n652));
  INV_X1    g466(.A(G472), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n538), .A2(new_n516), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n516), .A2(new_n522), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  AOI21_X1  g471(.A(G902), .B1(new_n657), .B2(new_n535), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n653), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n651), .A2(new_n652), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g474(.A(new_n645), .B(KEYINPUT39), .Z(new_n661));
  AND2_X1   g475(.A1(new_n309), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT40), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n381), .A2(new_n388), .ZN(new_n665));
  XOR2_X1   g479(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n666));
  XNOR2_X1  g480(.A(new_n665), .B(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n311), .ZN(new_n668));
  INV_X1    g482(.A(new_n491), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n626), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n639), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n664), .B(new_n672), .C1(new_n663), .C2(new_n662), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G143), .ZN(G45));
  INV_X1    g488(.A(KEYINPUT100), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n605), .A2(new_n491), .A3(new_n646), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n675), .B1(new_n648), .B2(new_n676), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n549), .A2(new_n309), .A3(new_n638), .ZN(new_n678));
  INV_X1    g492(.A(new_n676), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(KEYINPUT100), .A3(new_n611), .A4(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G146), .ZN(G48));
  OR2_X1    g496(.A1(new_n295), .A2(new_n190), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n297), .A2(new_n302), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n293), .B1(new_n305), .B2(new_n292), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n190), .B(new_n191), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n683), .A2(new_n188), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n688), .A2(new_n549), .A3(new_n584), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n690), .A2(KEYINPUT101), .A3(new_n611), .A4(new_n606), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n692), .B1(new_n612), .B2(new_n689), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT41), .B(G113), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G15));
  NAND4_X1  g510(.A1(new_n586), .A2(new_n627), .A3(new_n630), .A4(new_n688), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G116), .ZN(G18));
  NAND2_X1  g512(.A1(new_n611), .A2(new_n688), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n549), .A2(new_n492), .A3(new_n638), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(new_n317), .ZN(G21));
  INV_X1    g516(.A(KEYINPUT102), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n613), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n547), .A2(new_n191), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(KEYINPUT102), .A3(G472), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n536), .A2(new_n516), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n526), .A2(new_n523), .A3(new_n707), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n704), .A2(new_n706), .B1(new_n531), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n584), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n611), .A2(new_n688), .A3(new_n628), .A4(new_n670), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n392), .ZN(G24));
  NOR2_X1   g527(.A1(new_n699), .A2(new_n676), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT103), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n715), .B1(new_n709), .B2(new_n638), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n708), .A2(new_n531), .ZN(new_n717));
  AOI21_X1  g531(.A(KEYINPUT102), .B1(new_n705), .B2(G472), .ZN(new_n718));
  AOI211_X1 g532(.A(new_n703), .B(new_n653), .C1(new_n547), .C2(new_n191), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n638), .B(new_n717), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n720), .A2(KEYINPUT103), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n714), .B1(new_n716), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G125), .ZN(G27));
  NAND2_X1  g537(.A1(new_n543), .A2(new_n548), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(KEYINPUT106), .B2(new_n533), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n533), .A2(KEYINPUT106), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n583), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n303), .A2(G469), .A3(new_n306), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n189), .B1(new_n296), .B2(new_n728), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n381), .A2(new_n668), .A3(new_n388), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT104), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n192), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n686), .A2(new_n733), .A3(new_n728), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n188), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n381), .A2(new_n668), .A3(new_n388), .ZN(new_n736));
  OAI21_X1  g550(.A(KEYINPUT104), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n676), .B1(new_n732), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n727), .A2(KEYINPUT42), .A3(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n738), .A2(KEYINPUT105), .A3(new_n586), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT42), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(KEYINPUT105), .B1(new_n738), .B2(new_n586), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n739), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n744), .B(G131), .ZN(G33));
  NOR2_X1   g559(.A1(new_n647), .A2(new_n585), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n732), .A2(new_n737), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  AOI21_X1  g563(.A(KEYINPUT45), .B1(new_n300), .B2(new_n307), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n303), .A2(KEYINPUT45), .A3(new_n306), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(G469), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n733), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT46), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n753), .A2(new_n754), .B1(new_n190), .B2(new_n295), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n189), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n661), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT107), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n758), .B(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n605), .A2(new_n669), .ZN(new_n762));
  XOR2_X1   g576(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n763));
  NAND3_X1  g577(.A1(new_n762), .A2(KEYINPUT109), .A3(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n605), .A2(KEYINPUT43), .A3(new_n669), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(KEYINPUT109), .B1(new_n762), .B2(new_n763), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n761), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n767), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n769), .A2(KEYINPUT110), .A3(new_n765), .A4(new_n764), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n616), .A2(new_n639), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n768), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n760), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n768), .A2(new_n770), .A3(KEYINPUT44), .A4(new_n771), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n730), .B1(new_n776), .B2(KEYINPUT111), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT112), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(KEYINPUT111), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n778), .A2(new_n779), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n780), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT112), .B1(new_n782), .B2(new_n777), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n775), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(new_n236), .ZN(G39));
  NOR4_X1   g599(.A1(new_n676), .A2(new_n549), .A3(new_n584), .A4(new_n736), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT113), .Z(new_n787));
  XNOR2_X1  g601(.A(new_n757), .B(KEYINPUT47), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G140), .ZN(G42));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n791));
  INV_X1    g605(.A(new_n748), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT105), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n731), .B1(new_n729), .B2(new_n730), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n735), .A2(new_n736), .A3(KEYINPUT104), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n679), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n793), .B1(new_n796), .B2(new_n585), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n741), .A3(new_n740), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n792), .B1(new_n798), .B2(new_n739), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n389), .A2(new_n628), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n669), .A2(new_n625), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n801), .B(KEYINPUT116), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n621), .A2(new_n800), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n588), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n697), .A2(new_n641), .ZN(new_n805));
  OAI22_X1  g619(.A1(new_n710), .A2(new_n711), .B1(new_n699), .B2(new_n700), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n804), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT33), .B1(new_n427), .B2(new_n428), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n428), .A2(KEYINPUT94), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n809), .A2(KEYINPUT33), .A3(new_n593), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n426), .B(new_n594), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n808), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n603), .B1(new_n812), .B2(new_n599), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n604), .A2(new_n602), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n491), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(KEYINPUT114), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT114), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n605), .A2(new_n817), .A3(new_n491), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n800), .A3(new_n818), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n617), .B1(new_n819), .B2(KEYINPUT115), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT115), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n816), .A2(new_n800), .A3(new_n821), .A4(new_n818), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n693), .A2(new_n691), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n709), .A2(new_n715), .A3(new_n638), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n720), .A2(KEYINPUT103), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n626), .A2(new_n646), .ZN(new_n827));
  NOR4_X1   g641(.A1(new_n623), .A2(new_n827), .A3(new_n736), .A4(new_n624), .ZN(new_n828));
  AOI22_X1  g642(.A1(new_n826), .A2(new_n738), .B1(new_n678), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n799), .A2(new_n807), .A3(new_n823), .A4(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n649), .ZN(new_n831));
  AND2_X1   g645(.A1(new_n611), .A2(new_n670), .ZN(new_n832));
  INV_X1    g646(.A(new_n660), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n638), .A2(new_n735), .A3(new_n645), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n681), .A2(new_n722), .A3(new_n831), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT52), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n649), .B1(new_n826), .B2(new_n714), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n838), .A2(new_n839), .A3(new_n681), .A4(new_n835), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n791), .B1(new_n830), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n842), .A2(KEYINPUT119), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n837), .A2(new_n840), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n805), .A2(new_n806), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n803), .A2(new_n588), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n823), .A2(new_n845), .A3(new_n846), .A4(new_n829), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n744), .A2(new_n748), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n838), .A2(new_n839), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n844), .A2(new_n849), .A3(KEYINPUT53), .A4(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n852), .B(new_n791), .C1(new_n830), .C2(new_n841), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n843), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n854), .A2(KEYINPUT54), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n830), .A2(KEYINPUT117), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n830), .A2(KEYINPUT117), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n856), .A2(new_n857), .A3(new_n850), .A4(new_n844), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n846), .A2(new_n823), .A3(new_n845), .A4(new_n829), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n860), .A2(new_n799), .A3(new_n840), .A4(new_n837), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n859), .B1(new_n861), .B2(new_n791), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n844), .A2(new_n849), .A3(KEYINPUT118), .A4(KEYINPUT53), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n858), .A2(new_n791), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT54), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n855), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT51), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n766), .A2(new_n767), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n868), .A2(new_n441), .A3(new_n710), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n311), .A3(new_n667), .A4(new_n688), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT50), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(KEYINPUT120), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n871), .A2(KEYINPUT120), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n870), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n683), .A2(new_n686), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n875), .A2(new_n188), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n869), .B(new_n730), .C1(new_n788), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n687), .A2(new_n736), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n660), .A2(new_n584), .A3(new_n440), .A4(new_n879), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT121), .Z(new_n881));
  NOR2_X1   g695(.A1(new_n605), .A2(new_n491), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n868), .A2(new_n441), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n884), .A2(new_n826), .A3(new_n879), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n883), .B(new_n885), .C1(new_n872), .C2(new_n870), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n867), .B1(new_n878), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n884), .A2(new_n727), .A3(new_n879), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT48), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n869), .A2(new_n611), .A3(new_n688), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n881), .A2(new_n491), .A3(new_n605), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n891), .A2(G952), .A3(new_n193), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n887), .A2(new_n889), .A3(new_n890), .A4(new_n892), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n878), .A2(new_n886), .A3(new_n867), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI22_X1  g709(.A1(new_n866), .A2(new_n895), .B1(G952), .B2(G953), .ZN(new_n896));
  NOR3_X1   g710(.A1(new_n491), .A2(new_n311), .A3(new_n189), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n584), .B(new_n897), .C1(KEYINPUT49), .C2(new_n875), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(KEYINPUT49), .B2(new_n875), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n899), .A2(new_n605), .A3(new_n667), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n896), .B1(new_n833), .B2(new_n900), .ZN(G75));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n851), .A2(new_n853), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n852), .B1(new_n861), .B2(new_n791), .ZN(new_n904));
  OAI21_X1  g718(.A(G902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(G210), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n902), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n345), .A2(new_n356), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n354), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT55), .Z(new_n910));
  NAND2_X1  g724(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n197), .A2(G952), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT122), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n905), .A2(new_n915), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n854), .A2(KEYINPUT122), .A3(G902), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n916), .A2(new_n917), .A3(new_n313), .A4(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n910), .A2(KEYINPUT56), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n916), .A2(new_n313), .A3(new_n918), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT123), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n914), .B1(new_n921), .B2(new_n923), .ZN(G51));
  XNOR2_X1  g738(.A(new_n854), .B(new_n865), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n192), .B(KEYINPUT57), .Z(new_n926));
  OAI22_X1  g740(.A1(new_n925), .A2(new_n926), .B1(new_n685), .B2(new_n684), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n750), .A2(new_n752), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n916), .A2(new_n928), .A3(new_n918), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n912), .B1(new_n927), .B2(new_n929), .ZN(G54));
  AND2_X1   g744(.A1(KEYINPUT58), .A2(G475), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n916), .A2(new_n918), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n480), .A3(new_n473), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n916), .A2(new_n481), .A3(new_n918), .A4(new_n931), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n933), .A2(new_n913), .A3(new_n934), .ZN(G60));
  NAND2_X1  g749(.A1(G478), .A2(G902), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(KEYINPUT59), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n812), .B1(new_n866), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n812), .A2(new_n937), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n913), .B1(new_n925), .B2(new_n939), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n938), .A2(new_n940), .ZN(G63));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT60), .Z(new_n943));
  OAI211_X1 g757(.A(new_n636), .B(new_n943), .C1(new_n903), .C2(new_n904), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(KEYINPUT124), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT124), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n854), .A2(new_n946), .A3(new_n636), .A4(new_n943), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n577), .B1(new_n854), .B2(new_n943), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n949), .A2(new_n912), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT61), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n948), .A2(new_n950), .A3(KEYINPUT61), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(G66));
  INV_X1    g769(.A(new_n438), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n193), .B1(new_n956), .B2(G224), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n807), .A2(new_n823), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n957), .B1(new_n958), .B2(new_n197), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n908), .B1(G898), .B2(new_n197), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT125), .Z(new_n961));
  XNOR2_X1  g775(.A(new_n959), .B(new_n961), .ZN(G69));
  AOI21_X1  g776(.A(new_n197), .B1(G227), .B2(G900), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n519), .B1(new_n510), .B2(KEYINPUT30), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n464), .A2(new_n465), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n964), .B(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n966), .B1(new_n644), .B2(new_n197), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n848), .A2(KEYINPUT127), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n848), .A2(KEYINPUT127), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n760), .A2(new_n727), .A3(new_n832), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n968), .A2(new_n789), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n784), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n838), .A2(new_n681), .ZN(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n972), .A2(KEYINPUT126), .A3(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n976), .B1(new_n784), .B2(new_n973), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n971), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n967), .B1(new_n978), .B2(new_n197), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n974), .A2(new_n673), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n802), .B1(new_n816), .B2(new_n818), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n586), .A2(new_n662), .A3(new_n730), .ZN(new_n984));
  OR2_X1    g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n982), .A2(new_n789), .A3(new_n985), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n784), .A2(new_n981), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n987), .A2(new_n435), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n988), .A2(new_n966), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n963), .B1(new_n979), .B2(new_n989), .ZN(new_n990));
  OR2_X1    g804(.A1(new_n988), .A2(new_n966), .ZN(new_n991));
  INV_X1    g805(.A(new_n963), .ZN(new_n992));
  AOI211_X1 g806(.A(new_n435), .B(new_n971), .C1(new_n975), .C2(new_n977), .ZN(new_n993));
  OAI211_X1 g807(.A(new_n991), .B(new_n992), .C1(new_n993), .C2(new_n967), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n990), .A2(new_n994), .ZN(G72));
  NAND2_X1  g809(.A1(new_n657), .A2(new_n520), .ZN(new_n996));
  INV_X1    g810(.A(new_n958), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n978), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(G472), .A2(G902), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT63), .Z(new_n1000));
  AOI21_X1  g814(.A(new_n996), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  INV_X1    g815(.A(new_n525), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1000), .B1(new_n539), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1000), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n1004), .B1(new_n987), .B2(new_n997), .ZN(new_n1005));
  OAI221_X1 g819(.A(new_n913), .B1(new_n864), .B2(new_n1003), .C1(new_n1005), .C2(new_n655), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n1001), .A2(new_n1006), .ZN(G57));
endmodule


