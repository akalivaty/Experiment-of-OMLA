//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n821,
    new_n822, new_n824, new_n825, new_n826, new_n827, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(KEYINPUT77), .B(KEYINPUT30), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G226gat), .ZN(new_n208));
  INV_X1    g007(.A(G233gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT24), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(G183gat), .A3(G190gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(G183gat), .B(G190gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(new_n212), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n216));
  NAND2_X1  g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(G169gat), .ZN(new_n218));
  INV_X1    g017(.A(G176gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT23), .ZN(new_n220));
  OAI22_X1  g019(.A1(KEYINPUT67), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n221));
  AND2_X1   g020(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n217), .B(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT68), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT66), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n226), .B(new_n213), .C1(new_n214), .C2(new_n212), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n216), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT25), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n215), .A2(KEYINPUT25), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n223), .B1(new_n224), .B2(new_n229), .ZN(new_n231));
  AOI22_X1  g030(.A1(new_n228), .A2(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT27), .B(G183gat), .ZN(new_n233));
  INV_X1    g032(.A(G190gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT28), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(G183gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(new_n234), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT26), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n217), .A2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  AOI211_X1 g042(.A(new_n239), .B(new_n243), .C1(KEYINPUT26), .C2(new_n242), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n237), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n232), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n211), .B1(new_n246), .B2(KEYINPUT29), .ZN(new_n247));
  XNOR2_X1  g046(.A(G197gat), .B(G204gat), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT22), .ZN(new_n249));
  INV_X1    g048(.A(G211gat), .ZN(new_n250));
  INV_X1    g049(.A(G218gat), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G211gat), .B(G218gat), .ZN(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n254), .A2(new_n248), .A3(new_n252), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT75), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n256), .A2(KEYINPUT75), .A3(new_n257), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT76), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n264), .B(new_n210), .C1(new_n232), .C2(new_n245), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n237), .A2(new_n244), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n212), .A2(G183gat), .A3(G190gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n238), .A2(G190gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n234), .A2(G183gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(new_n268), .B1(new_n271), .B2(KEYINPUT24), .ZN(new_n272));
  AOI22_X1  g071(.A1(new_n272), .A2(new_n226), .B1(new_n223), .B2(new_n224), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT25), .B1(new_n273), .B2(new_n216), .ZN(new_n274));
  AND2_X1   g073(.A1(new_n231), .A2(new_n230), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n267), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n264), .B1(new_n276), .B2(new_n210), .ZN(new_n277));
  OAI211_X1 g076(.A(new_n247), .B(new_n263), .C1(new_n266), .C2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT29), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n210), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n228), .A2(new_n229), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n231), .A2(new_n230), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n211), .B1(new_n283), .B2(new_n267), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n262), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  AOI211_X1 g084(.A(new_n205), .B(new_n207), .C1(new_n278), .C2(new_n285), .ZN(new_n286));
  AND2_X1   g085(.A1(new_n278), .A2(new_n285), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n205), .ZN(new_n288));
  NAND2_X1  g087(.A1(KEYINPUT77), .A2(KEYINPUT30), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n278), .A2(new_n285), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(new_n204), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n286), .B1(new_n288), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n294));
  INV_X1    g093(.A(G113gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n294), .B1(new_n295), .B2(G120gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(G120gat), .ZN(new_n297));
  INV_X1    g096(.A(G120gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n298), .A2(KEYINPUT71), .A3(G113gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n296), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  OR2_X1    g099(.A1(new_n300), .A2(KEYINPUT72), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(KEYINPUT72), .ZN(new_n302));
  XNOR2_X1  g101(.A(G127gat), .B(G134gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT1), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(new_n302), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT70), .ZN(new_n308));
  INV_X1    g107(.A(G134gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G127gat), .ZN(new_n310));
  INV_X1    g109(.A(G127gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G134gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT69), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT69), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n303), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n295), .A2(G120gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n298), .A2(G113gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n304), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n308), .B1(new_n317), .B2(new_n320), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n310), .A2(new_n312), .A3(new_n315), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n315), .B1(new_n310), .B2(new_n312), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n308), .B(new_n320), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n307), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT78), .ZN(new_n327));
  INV_X1    g126(.A(G148gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n327), .B1(new_n328), .B2(G141gat), .ZN(new_n329));
  INV_X1    g128(.A(G141gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n330), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n329), .B(new_n331), .C1(new_n330), .C2(G148gat), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT2), .ZN(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(new_n334), .B2(new_n335), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n332), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n328), .A2(G141gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n330), .A2(G148gat), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n333), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  XOR2_X1   g140(.A(G155gat), .B(G162gat), .Z(new_n342));
  NAND2_X1  g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  OR2_X1    g143(.A1(new_n344), .A2(KEYINPUT3), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n326), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(KEYINPUT5), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n338), .A2(new_n343), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n307), .B(new_n352), .C1(new_n321), .C2(new_n325), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT80), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n356), .A2(KEYINPUT70), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n324), .ZN(new_n358));
  NAND4_X1  g157(.A1(new_n358), .A2(KEYINPUT80), .A3(new_n307), .A4(new_n352), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n351), .B1(new_n355), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n338), .A2(new_n343), .A3(KEYINPUT79), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g161(.A(KEYINPUT79), .B1(new_n338), .B2(new_n343), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n305), .B1(new_n300), .B2(KEYINPUT72), .ZN(new_n365));
  AOI22_X1  g164(.A1(new_n357), .A2(new_n324), .B1(new_n301), .B2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n366), .A3(new_n351), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n350), .B1(new_n360), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G1gat), .B(G29gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n370), .B(KEYINPUT0), .ZN(new_n371));
  XNOR2_X1  g170(.A(G57gat), .B(G85gat), .ZN(new_n372));
  XOR2_X1   g171(.A(new_n371), .B(new_n372), .Z(new_n373));
  OAI21_X1  g172(.A(KEYINPUT81), .B1(new_n366), .B2(new_n352), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n326), .A2(new_n375), .A3(new_n344), .ZN(new_n376));
  AOI22_X1  g175(.A1(new_n374), .A2(new_n376), .B1(new_n355), .B2(new_n359), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT5), .B1(new_n377), .B2(new_n348), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT4), .B1(new_n355), .B2(new_n359), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n364), .A2(new_n366), .A3(KEYINPUT4), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(new_n347), .A3(new_n348), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n369), .B(new_n373), .C1(new_n378), .C2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT5), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n374), .A2(new_n376), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n355), .A2(new_n359), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(new_n348), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n385), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  OR2_X1    g189(.A1(new_n379), .A2(new_n381), .ZN(new_n391));
  OR2_X1    g190(.A1(new_n360), .A2(new_n368), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n390), .A2(new_n391), .B1(new_n392), .B2(new_n350), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n383), .B(new_n384), .C1(new_n393), .C2(new_n373), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n369), .B1(new_n378), .B2(new_n382), .ZN(new_n395));
  INV_X1    g194(.A(new_n373), .ZN(new_n396));
  INV_X1    g195(.A(new_n384), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n293), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g199(.A(KEYINPUT31), .B(G50gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n279), .B1(new_n344), .B2(KEYINPUT3), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(new_n261), .A3(new_n260), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT29), .B1(new_n256), .B2(new_n257), .ZN(new_n404));
  OAI22_X1  g203(.A1(new_n362), .A2(new_n363), .B1(new_n404), .B2(KEYINPUT3), .ZN(new_n405));
  NAND2_X1  g204(.A1(G228gat), .A2(G233gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n403), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n344), .B1(new_n404), .B2(KEYINPUT3), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n406), .B1(new_n403), .B2(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n401), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n410), .ZN(new_n412));
  INV_X1    g211(.A(new_n401), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n407), .A3(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G78gat), .B(G106gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(G22gat), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n411), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n416), .B1(new_n411), .B2(new_n414), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n400), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT36), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n283), .A2(new_n326), .A3(new_n267), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n366), .B1(new_n232), .B2(new_n245), .ZN(new_n424));
  NAND2_X1  g223(.A1(G227gat), .A2(G233gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT64), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n426), .B(KEYINPUT65), .ZN(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n423), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT32), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT33), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(G15gat), .B(G43gat), .Z(new_n433));
  XNOR2_X1  g232(.A(G71gat), .B(G99gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n430), .A2(new_n432), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n435), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n429), .B(KEYINPUT32), .C1(new_n431), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  OR2_X1    g240(.A1(new_n428), .A2(KEYINPUT34), .ZN(new_n442));
  OR2_X1    g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(KEYINPUT73), .B(KEYINPUT34), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n426), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n445), .B1(new_n441), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n443), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n439), .A2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n436), .A2(new_n443), .A3(new_n447), .A4(new_n438), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n422), .B1(new_n452), .B2(KEYINPUT74), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT74), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n454), .A3(KEYINPUT36), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n421), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n263), .B1(new_n280), .B2(new_n284), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n247), .B(new_n262), .C1(new_n266), .C2(new_n277), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n457), .A2(new_n458), .ZN(new_n462));
  OAI21_X1  g261(.A(KEYINPUT37), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT38), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n205), .A2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT37), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n290), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n290), .A2(new_n204), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(new_n394), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n398), .A2(KEYINPUT84), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT84), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n395), .A2(new_n472), .A3(new_n396), .A4(new_n397), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n287), .A2(KEYINPUT37), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n204), .B1(new_n290), .B2(new_n466), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n464), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n470), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT40), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n347), .B1(new_n360), .B2(new_n368), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT39), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n389), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n373), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n386), .A2(new_n387), .A3(new_n348), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT39), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n485), .B1(new_n389), .B2(new_n480), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n479), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n480), .A2(new_n389), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n488), .A2(KEYINPUT39), .A3(new_n484), .ZN(new_n489));
  NAND4_X1  g288(.A1(new_n489), .A2(KEYINPUT40), .A3(new_n373), .A4(new_n482), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n395), .A2(new_n396), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n487), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n419), .B1(new_n293), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT85), .B1(new_n478), .B2(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n471), .A2(new_n473), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n394), .A2(new_n469), .ZN(new_n496));
  INV_X1    g295(.A(new_n477), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n495), .A2(new_n496), .A3(new_n497), .A4(new_n468), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n487), .A2(new_n491), .A3(new_n490), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n420), .B1(new_n499), .B2(new_n292), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT85), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n456), .B1(new_n494), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n449), .A2(new_n419), .A3(new_n450), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n504), .A2(new_n292), .ZN(new_n505));
  XOR2_X1   g304(.A(KEYINPUT86), .B(KEYINPUT35), .Z(new_n506));
  NAND3_X1  g305(.A1(new_n471), .A2(new_n394), .A3(new_n473), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n505), .A2(KEYINPUT87), .A3(new_n506), .A4(new_n507), .ZN(new_n511));
  OAI21_X1  g310(.A(KEYINPUT35), .B1(new_n400), .B2(new_n504), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n503), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G15gat), .B(G22gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT16), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(G1gat), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n517), .B1(G1gat), .B2(new_n515), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(G8gat), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G36gat), .ZN(new_n521));
  AND2_X1   g320(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n521), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G29gat), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n528));
  XNOR2_X1  g327(.A(G43gat), .B(G50gat), .ZN(new_n529));
  OR2_X1    g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n527), .A2(KEYINPUT15), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n528), .A2(new_n529), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n533), .A2(KEYINPUT88), .A3(KEYINPUT17), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT17), .B1(new_n533), .B2(KEYINPUT88), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n520), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(G229gat), .A2(G233gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n533), .A2(new_n519), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n536), .A2(KEYINPUT18), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  OR3_X1    g338(.A1(new_n533), .A2(new_n519), .A3(KEYINPUT90), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT90), .B1(new_n533), .B2(new_n519), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(new_n537), .B(KEYINPUT13), .Z(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n536), .A2(new_n537), .A3(new_n538), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT18), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n539), .A2(new_n544), .A3(KEYINPUT89), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G197gat), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT11), .B(G169gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT12), .Z(new_n555));
  NAND3_X1  g354(.A1(new_n549), .A2(new_n550), .A3(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(new_n555), .ZN(new_n557));
  OAI211_X1 g356(.A(new_n545), .B(new_n548), .C1(KEYINPUT89), .C2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  AND2_X1   g358(.A1(new_n514), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(G232gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n561), .A2(new_n209), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n562), .A2(KEYINPUT41), .ZN(new_n563));
  XNOR2_X1  g362(.A(G134gat), .B(G162gat), .ZN(new_n564));
  XOR2_X1   g363(.A(new_n563), .B(new_n564), .Z(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  INV_X1    g367(.A(G92gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT95), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT94), .B(KEYINPUT7), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n568), .A2(new_n569), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G99gat), .B(G106gat), .Z(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n576), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n571), .A2(new_n574), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n533), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n562), .A2(KEYINPUT41), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n580), .B1(new_n534), .B2(new_n535), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT96), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g386(.A(KEYINPUT96), .B(new_n580), .C1(new_n534), .C2(new_n535), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G190gat), .B(G218gat), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(KEYINPUT93), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n589), .A2(new_n590), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n566), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G71gat), .A2(G78gat), .ZN(new_n595));
  OR2_X1    g394(.A1(G71gat), .A2(G78gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT9), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G57gat), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(G64gat), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(G64gat), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n600), .B1(new_n601), .B2(KEYINPUT91), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT91), .ZN(new_n603));
  NOR3_X1   g402(.A1(new_n603), .A2(new_n599), .A3(G64gat), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n598), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(G64gat), .ZN(new_n606));
  NOR2_X1   g405(.A1(new_n606), .A2(G57gat), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT9), .B1(new_n601), .B2(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n608), .A2(new_n595), .A3(new_n596), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT21), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(G231gat), .A2(G233gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G127gat), .B(G155gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT92), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n614), .B(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G183gat), .B(G211gat), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n520), .B1(new_n611), .B2(new_n610), .ZN(new_n620));
  XOR2_X1   g419(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  OR2_X1    g423(.A1(new_n617), .A2(new_n618), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n617), .A2(new_n618), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n625), .A2(new_n622), .A3(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n589), .A2(new_n590), .ZN(new_n629));
  NAND4_X1  g428(.A1(new_n629), .A2(KEYINPUT93), .A3(new_n591), .A4(new_n565), .ZN(new_n630));
  XNOR2_X1  g429(.A(G120gat), .B(G148gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(G176gat), .B(G204gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT10), .ZN(new_n635));
  NOR3_X1   g434(.A1(new_n580), .A2(new_n635), .A3(new_n610), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n575), .A2(KEYINPUT97), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n576), .ZN(new_n638));
  INV_X1    g437(.A(new_n610), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n637), .A2(new_n576), .ZN(new_n641));
  OAI22_X1  g440(.A1(new_n640), .A2(new_n641), .B1(new_n580), .B2(new_n639), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n636), .B1(new_n642), .B2(new_n635), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n644), .B(KEYINPUT98), .Z(new_n645));
  NOR2_X1   g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n640), .A2(new_n641), .ZN(new_n647));
  INV_X1    g446(.A(new_n644), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n581), .A2(new_n610), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n634), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  OAI211_X1 g451(.A(new_n650), .B(new_n633), .C1(new_n643), .C2(new_n648), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n594), .A2(new_n628), .A3(new_n630), .A4(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n560), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n399), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G1gat), .ZN(G1324gat));
  NOR2_X1   g461(.A1(new_n658), .A2(new_n293), .ZN(new_n663));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(G8gat), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n665), .B1(new_n666), .B2(new_n663), .ZN(new_n667));
  MUX2_X1   g466(.A(new_n665), .B(new_n667), .S(KEYINPUT42), .Z(G1325gat));
  AOI21_X1  g467(.A(G15gat), .B1(new_n659), .B2(new_n452), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n453), .A2(new_n455), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(G15gat), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(KEYINPUT99), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n669), .B1(new_n659), .B2(new_n672), .ZN(G1326gat));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n419), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT43), .B(G22gat), .Z(new_n675));
  XNOR2_X1  g474(.A(new_n674), .B(new_n675), .ZN(G1327gat));
  NAND2_X1  g475(.A1(new_n594), .A2(new_n630), .ZN(new_n677));
  INV_X1    g476(.A(new_n628), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(new_n678), .A3(new_n655), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT100), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n560), .A2(new_n680), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n681), .A2(G29gat), .A3(new_n399), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT45), .Z(new_n683));
  OAI21_X1  g482(.A(new_n677), .B1(new_n503), .B2(new_n513), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI211_X1 g485(.A(KEYINPUT44), .B(new_n677), .C1(new_n503), .C2(new_n513), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n654), .B(KEYINPUT101), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n559), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n689), .A2(new_n690), .A3(new_n628), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n686), .A2(new_n687), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT102), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n686), .A2(KEYINPUT102), .A3(new_n687), .A4(new_n691), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n694), .A2(new_n660), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n683), .B1(new_n525), .B2(new_n696), .ZN(G1328gat));
  NAND4_X1  g496(.A1(new_n560), .A2(new_n521), .A3(new_n292), .A4(new_n680), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(KEYINPUT46), .ZN(new_n699));
  OR2_X1    g498(.A1(new_n698), .A2(KEYINPUT46), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n694), .A2(new_n292), .A3(new_n695), .ZN(new_n701));
  OAI211_X1 g500(.A(new_n699), .B(new_n700), .C1(new_n701), .C2(new_n521), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1329gat));
  NOR3_X1   g503(.A1(new_n681), .A2(G43gat), .A3(new_n451), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n694), .A2(new_n670), .A3(new_n695), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(G43gat), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT47), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  INV_X1    g508(.A(G43gat), .ZN(new_n710));
  INV_X1    g509(.A(new_n692), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n710), .B1(new_n711), .B2(new_n670), .ZN(new_n712));
  OAI22_X1  g511(.A1(KEYINPUT47), .A2(new_n707), .B1(new_n709), .B2(new_n712), .ZN(G1330gat));
  NOR3_X1   g512(.A1(new_n681), .A2(G50gat), .A3(new_n419), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT48), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G50gat), .B1(new_n692), .B2(new_n419), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n694), .A2(new_n420), .A3(new_n695), .ZN(new_n719));
  AND3_X1   g518(.A1(new_n719), .A2(KEYINPUT104), .A3(G50gat), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT104), .B1(new_n719), .B2(G50gat), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n720), .A2(new_n721), .A3(new_n714), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n718), .B1(new_n722), .B2(KEYINPUT48), .ZN(G1331gat));
  NOR4_X1   g522(.A1(new_n688), .A2(new_n677), .A3(new_n678), .A4(new_n559), .ZN(new_n724));
  AND2_X1   g523(.A1(new_n514), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n660), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g526(.A1(new_n725), .A2(new_n292), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n728), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT49), .B(G64gat), .Z(new_n730));
  OAI21_X1  g529(.A(new_n729), .B1(new_n728), .B2(new_n730), .ZN(G1333gat));
  NAND2_X1  g530(.A1(new_n725), .A2(new_n670), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n451), .A2(G71gat), .ZN(new_n733));
  AOI22_X1  g532(.A1(new_n732), .A2(G71gat), .B1(new_n725), .B2(new_n733), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g534(.A1(new_n725), .A2(new_n420), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(G78gat), .ZN(G1335gat));
  AND2_X1   g536(.A1(new_n686), .A2(new_n687), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n559), .A2(new_n628), .A3(new_n655), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(G85gat), .B1(new_n740), .B2(new_n399), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n559), .A2(new_n628), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n514), .A2(new_n677), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g544(.A1(new_n514), .A2(KEYINPUT51), .A3(new_n677), .A4(new_n742), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(KEYINPUT105), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT105), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n743), .A2(new_n748), .A3(new_n744), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n660), .A2(new_n568), .A3(new_n654), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n741), .B1(new_n750), .B2(new_n751), .ZN(G1336gat));
  NAND3_X1  g551(.A1(new_n738), .A2(new_n292), .A3(new_n739), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n753), .A2(new_n754), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n755), .A2(new_n756), .A3(new_n569), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n688), .A2(G92gat), .A3(new_n293), .ZN(new_n759));
  INV_X1    g558(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n750), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n762));
  AOI22_X1  g561(.A1(new_n753), .A2(G92gat), .B1(new_n762), .B2(new_n759), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n757), .A2(new_n761), .B1(new_n758), .B2(new_n763), .ZN(G1337gat));
  AOI21_X1  g563(.A(new_n740), .B1(new_n453), .B2(new_n455), .ZN(new_n765));
  XNOR2_X1  g564(.A(KEYINPUT107), .B(G99gat), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n452), .A2(new_n654), .A3(new_n766), .ZN(new_n767));
  OAI22_X1  g566(.A1(new_n765), .A2(new_n766), .B1(new_n750), .B2(new_n767), .ZN(G1338gat));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  OAI21_X1  g568(.A(G106gat), .B1(new_n740), .B2(new_n419), .ZN(new_n770));
  NOR3_X1   g569(.A1(new_n688), .A2(G106gat), .A3(new_n419), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n747), .A2(new_n749), .A3(new_n771), .ZN(new_n772));
  AND2_X1   g571(.A1(new_n772), .A2(KEYINPUT108), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(KEYINPUT108), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n769), .B(new_n770), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n762), .A2(new_n771), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n770), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT53), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n775), .A2(new_n778), .ZN(G1339gat));
  INV_X1    g578(.A(new_n677), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n537), .B1(new_n536), .B2(new_n538), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT110), .ZN(new_n782));
  OAI22_X1  g581(.A1(new_n781), .A2(new_n782), .B1(new_n543), .B2(new_n542), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n554), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n545), .A2(new_n548), .A3(new_n557), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(new_n654), .ZN(new_n788));
  OAI21_X1  g587(.A(KEYINPUT54), .B1(new_n643), .B2(new_n648), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n643), .A2(new_n645), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(new_n792), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT109), .B1(new_n794), .B2(new_n789), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n646), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n634), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n796), .A2(KEYINPUT55), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n653), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n799), .B1(new_n793), .B2(new_n795), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n559), .B1(new_n803), .B2(KEYINPUT55), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n780), .B(new_n788), .C1(new_n802), .C2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n787), .B1(new_n803), .B2(KEYINPUT55), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n677), .B1(new_n802), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(new_n807), .A3(new_n678), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n808), .B1(new_n559), .B2(new_n656), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n809), .A2(new_n419), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n810), .A2(new_n660), .A3(new_n293), .A4(new_n452), .ZN(new_n811));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n690), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n809), .A2(new_n660), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n813), .A2(new_n292), .A3(new_n504), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(new_n295), .A3(new_n559), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n812), .A2(new_n815), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT111), .Z(G1340gat));
  NOR3_X1   g616(.A1(new_n811), .A2(new_n298), .A3(new_n688), .ZN(new_n818));
  AOI21_X1  g617(.A(G120gat), .B1(new_n814), .B2(new_n654), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n818), .A2(new_n819), .ZN(G1341gat));
  OAI21_X1  g619(.A(G127gat), .B1(new_n811), .B2(new_n678), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n814), .A2(new_n311), .A3(new_n628), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1342gat));
  NAND2_X1  g622(.A1(new_n293), .A2(new_n309), .ZN(new_n824));
  NOR4_X1   g623(.A1(new_n813), .A2(new_n504), .A3(new_n780), .A4(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT56), .ZN(new_n826));
  OAI21_X1  g625(.A(G134gat), .B1(new_n811), .B2(new_n780), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(G1343gat));
  INV_X1    g627(.A(new_n813), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n670), .A2(new_n292), .A3(new_n419), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n831), .A2(G141gat), .A3(new_n690), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n809), .A2(new_n420), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n833), .A2(KEYINPUT57), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n670), .A2(new_n399), .A3(new_n292), .ZN(new_n835));
  XOR2_X1   g634(.A(KEYINPUT112), .B(KEYINPUT57), .Z(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n834), .A2(new_n835), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT113), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT113), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n834), .A2(new_n841), .A3(new_n835), .A4(new_n838), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n559), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n832), .B1(new_n843), .B2(G141gat), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  XNOR2_X1  g644(.A(KEYINPUT114), .B(KEYINPUT58), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n832), .A2(new_n846), .ZN(new_n847));
  OAI21_X1  g646(.A(G141gat), .B1(new_n839), .B2(new_n690), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT115), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n847), .B2(new_n848), .ZN(new_n851));
  OAI22_X1  g650(.A1(new_n844), .A2(new_n845), .B1(new_n850), .B2(new_n851), .ZN(G1344gat));
  INV_X1    g651(.A(new_n831), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n853), .A2(new_n328), .A3(new_n654), .ZN(new_n854));
  OR2_X1    g653(.A1(new_n328), .A2(KEYINPUT59), .ZN(new_n855));
  AND2_X1   g654(.A1(new_n840), .A2(new_n842), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n856), .B2(new_n654), .ZN(new_n857));
  XNOR2_X1  g656(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n858));
  OR3_X1    g657(.A1(new_n656), .A2(KEYINPUT117), .A3(new_n559), .ZN(new_n859));
  OAI21_X1  g658(.A(KEYINPUT117), .B1(new_n656), .B2(new_n559), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n808), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n419), .B1(new_n862), .B2(KEYINPUT118), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT118), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n808), .A2(new_n861), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT57), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n809), .A2(new_n420), .A3(new_n837), .ZN(new_n867));
  INV_X1    g666(.A(new_n867), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n654), .B(new_n835), .C1(new_n866), .C2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n858), .B1(new_n869), .B2(G148gat), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n854), .B1(new_n857), .B2(new_n870), .ZN(G1345gat));
  AOI21_X1  g670(.A(G155gat), .B1(new_n853), .B2(new_n628), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n628), .A2(G155gat), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT119), .Z(new_n874));
  AOI21_X1  g673(.A(new_n872), .B1(new_n856), .B2(new_n874), .ZN(G1346gat));
  NAND3_X1  g674(.A1(new_n853), .A2(new_n335), .A3(new_n677), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n856), .A2(new_n677), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n876), .B1(new_n877), .B2(new_n335), .ZN(G1347gat));
  NAND2_X1  g677(.A1(new_n399), .A2(new_n292), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT120), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n451), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n810), .A2(new_n881), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(new_n218), .A3(new_n690), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n809), .A2(new_n399), .ZN(new_n884));
  AND4_X1   g683(.A1(new_n292), .A2(new_n884), .A3(new_n419), .A4(new_n452), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n559), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n883), .B1(new_n218), .B2(new_n886), .ZN(G1348gat));
  NAND3_X1  g686(.A1(new_n885), .A2(new_n219), .A3(new_n654), .ZN(new_n888));
  OAI21_X1  g687(.A(G176gat), .B1(new_n882), .B2(new_n688), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g689(.A(new_n890), .B(KEYINPUT121), .Z(G1349gat));
  NAND3_X1  g690(.A1(new_n885), .A2(new_n233), .A3(new_n628), .ZN(new_n892));
  OAI21_X1  g691(.A(G183gat), .B1(new_n882), .B2(new_n678), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g694(.A(G190gat), .B1(new_n882), .B2(new_n780), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT122), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n900), .B1(new_n897), .B2(new_n896), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n898), .A2(new_n899), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n234), .A3(new_n677), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(G1351gat));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n905), .B1(new_n866), .B2(new_n868), .ZN(new_n906));
  AND3_X1   g705(.A1(new_n808), .A2(new_n861), .A3(new_n864), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n864), .B1(new_n808), .B2(new_n861), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n907), .A2(new_n908), .A3(new_n419), .ZN(new_n909));
  OAI211_X1 g708(.A(KEYINPUT123), .B(new_n867), .C1(new_n909), .C2(KEYINPUT57), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n880), .A2(new_n670), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n906), .A2(new_n910), .A3(new_n559), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(G197gat), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n670), .A2(new_n293), .A3(new_n419), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n884), .A2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(G197gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n916), .A3(new_n559), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(KEYINPUT124), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n913), .A2(new_n920), .A3(new_n917), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n919), .A2(new_n921), .ZN(G1352gat));
  INV_X1    g721(.A(G204gat), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n915), .A2(new_n923), .A3(new_n654), .ZN(new_n924));
  XOR2_X1   g723(.A(KEYINPUT125), .B(KEYINPUT62), .Z(new_n925));
  XNOR2_X1  g724(.A(new_n924), .B(new_n925), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT126), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n906), .A2(new_n910), .A3(new_n911), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n928), .B2(new_n688), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(G204gat), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n928), .A2(new_n927), .A3(new_n688), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n926), .B1(new_n930), .B2(new_n931), .ZN(G1353gat));
  NAND3_X1  g731(.A1(new_n915), .A2(new_n250), .A3(new_n628), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n911), .A2(new_n628), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n934), .B(new_n936), .C1(new_n866), .C2(new_n868), .ZN(new_n937));
  AND2_X1   g736(.A1(new_n937), .A2(G211gat), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n936), .B1(new_n866), .B2(new_n868), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n939), .A2(KEYINPUT127), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n938), .A2(KEYINPUT63), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n938), .B2(new_n940), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n933), .B1(new_n941), .B2(new_n942), .ZN(G1354gat));
  NOR3_X1   g742(.A1(new_n928), .A2(new_n251), .A3(new_n780), .ZN(new_n944));
  AOI21_X1  g743(.A(G218gat), .B1(new_n915), .B2(new_n677), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n944), .A2(new_n945), .ZN(G1355gat));
endmodule


