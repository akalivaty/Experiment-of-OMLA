//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 0 0 1 1 1 1 1 1 1 0 1 0 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n756, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n805, new_n806, new_n807, new_n808, new_n809, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n187));
  INV_X1    g001(.A(G217), .ZN(new_n188));
  INV_X1    g002(.A(G902), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n188), .B1(G234), .B2(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(KEYINPUT75), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT75), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(G125), .A3(G140), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n192), .B1(new_n195), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NOR3_X1   g013(.A1(new_n194), .A2(KEYINPUT16), .A3(G140), .ZN(new_n200));
  OR3_X1    g014(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n199), .B1(new_n198), .B2(new_n200), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT74), .B1(new_n204), .B2(G128), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT23), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n204), .A2(G128), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT23), .ZN(new_n208));
  OAI211_X1 g022(.A(KEYINPUT74), .B(new_n208), .C1(new_n204), .C2(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  XOR2_X1   g024(.A(KEYINPUT24), .B(G110), .Z(new_n211));
  XNOR2_X1  g025(.A(G119), .B(G128), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI22_X1  g027(.A1(G110), .A2(new_n210), .B1(new_n213), .B2(KEYINPUT73), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n203), .A2(new_n214), .ZN(new_n215));
  OR2_X1    g029(.A1(new_n213), .A2(KEYINPUT73), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G137), .ZN(new_n218));
  INV_X1    g032(.A(G953), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT68), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT68), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G953), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(G221), .A3(G234), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT22), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n224), .A2(KEYINPUT22), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n218), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n227), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n229), .A2(G137), .A3(new_n225), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G110), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n206), .A2(new_n233), .A3(new_n207), .A4(new_n209), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT76), .ZN(new_n235));
  OR2_X1    g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n235), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n236), .B(new_n237), .C1(new_n212), .C2(new_n211), .ZN(new_n238));
  NOR3_X1   g052(.A1(new_n198), .A2(new_n199), .A3(new_n200), .ZN(new_n239));
  XNOR2_X1  g053(.A(G125), .B(G140), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n239), .B1(new_n199), .B2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n217), .A2(new_n232), .A3(new_n242), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n228), .A2(new_n230), .A3(KEYINPUT77), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT77), .B1(new_n228), .B2(new_n230), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n215), .A2(new_n216), .B1(new_n238), .B2(new_n241), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n243), .B(new_n189), .C1(new_n246), .C2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT25), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n217), .A2(new_n242), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n251), .B1(new_n244), .B2(new_n245), .ZN(new_n252));
  NAND4_X1  g066(.A1(new_n252), .A2(KEYINPUT25), .A3(new_n189), .A4(new_n243), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n191), .B1(new_n250), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n243), .ZN(new_n256));
  NOR3_X1   g070(.A1(new_n256), .A2(G902), .A3(new_n190), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n187), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  NOR3_X1   g073(.A1(new_n254), .A2(new_n257), .A3(KEYINPUT78), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT30), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n263));
  INV_X1    g077(.A(G143), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G146), .ZN(new_n265));
  AND2_X1   g079(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n266));
  NOR2_X1   g080(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n199), .A2(G143), .ZN(new_n269));
  AOI21_X1  g083(.A(G128), .B1(new_n269), .B2(new_n265), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n263), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OR2_X1    g085(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n272));
  NAND2_X1  g086(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n272), .A2(new_n264), .A3(G146), .A4(new_n273), .ZN(new_n274));
  XNOR2_X1  g088(.A(G143), .B(G146), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n274), .B(KEYINPUT66), .C1(G128), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n272), .A2(new_n273), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n275), .A3(G128), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n271), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G131), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT11), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(KEYINPUT64), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT64), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G134), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n283), .A2(new_n285), .A3(G137), .ZN(new_n286));
  NOR2_X1   g100(.A1(G134), .A2(G137), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n281), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT64), .B(G134), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n290), .A2(new_n281), .A3(new_n218), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n280), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n282), .A2(G137), .ZN(new_n293));
  INV_X1    g107(.A(new_n290), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n293), .B1(new_n294), .B2(G137), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G131), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n279), .A2(new_n292), .A3(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n275), .A2(KEYINPUT0), .A3(G128), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT0), .B(G128), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n298), .B1(new_n275), .B2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n290), .A2(new_n281), .A3(new_n218), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n287), .B1(new_n290), .B2(G137), .ZN(new_n302));
  OAI211_X1 g116(.A(G131), .B(new_n301), .C1(new_n302), .C2(new_n281), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n300), .B1(new_n292), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n262), .B1(new_n297), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n292), .A2(new_n303), .ZN(new_n306));
  INV_X1    g120(.A(new_n300), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n279), .A2(new_n292), .A3(new_n296), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n308), .A2(KEYINPUT30), .A3(new_n309), .ZN(new_n310));
  OR2_X1    g124(.A1(KEYINPUT2), .A2(G113), .ZN(new_n311));
  NAND2_X1  g125(.A1(KEYINPUT2), .A2(G113), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n204), .A2(G116), .ZN(new_n314));
  INV_X1    g128(.A(G116), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n317), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n311), .A2(new_n314), .A3(new_n316), .A4(new_n312), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n305), .A2(new_n310), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G237), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n223), .A2(G210), .A3(new_n322), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT27), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(KEYINPUT26), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT27), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n323), .B(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT26), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n325), .A2(new_n329), .A3(G101), .ZN(new_n330));
  AOI21_X1  g144(.A(G101), .B1(new_n325), .B2(new_n329), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT67), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n320), .B(new_n333), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n308), .A2(new_n309), .A3(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n321), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(KEYINPUT31), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT28), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n320), .B1(new_n297), .B2(new_n304), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n308), .A2(new_n334), .A3(KEYINPUT28), .A4(new_n309), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n332), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT31), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n321), .A2(new_n332), .A3(new_n345), .A4(new_n335), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n337), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(G472), .A2(G902), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT69), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n347), .A2(new_n351), .A3(new_n348), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n351), .B1(new_n347), .B2(new_n348), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n349), .A2(KEYINPUT69), .A3(new_n351), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT72), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT71), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n339), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n335), .A2(KEYINPUT71), .A3(new_n338), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n330), .A2(new_n331), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT70), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n320), .B(KEYINPUT67), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n297), .B2(new_n304), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n335), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n365), .B1(new_n368), .B2(KEYINPUT28), .ZN(new_n369));
  AOI211_X1 g183(.A(KEYINPUT70), .B(new_n338), .C1(new_n367), .C2(new_n335), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n362), .B(new_n364), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n358), .B1(new_n371), .B2(new_n189), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  OR2_X1    g187(.A1(new_n342), .A2(new_n343), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n321), .A2(new_n335), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n343), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n374), .A2(new_n363), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n371), .A2(new_n358), .A3(new_n189), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n373), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G472), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n261), .B1(new_n357), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G469), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n223), .A2(G227), .ZN(new_n383));
  XNOR2_X1  g197(.A(G110), .B(G140), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT80), .ZN(new_n386));
  INV_X1    g200(.A(G107), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(new_n387), .A3(G104), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n388), .A2(KEYINPUT3), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n387), .A2(G104), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n386), .A2(new_n392), .A3(new_n387), .A4(G104), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT81), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT81), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n389), .A2(new_n396), .A3(new_n391), .A4(new_n393), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(G101), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G101), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n389), .A2(new_n399), .A3(new_n391), .A4(new_n393), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(KEYINPUT4), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n300), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(G104), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(G107), .ZN(new_n407));
  OAI21_X1  g221(.A(G101), .B1(new_n390), .B2(new_n407), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n400), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n279), .A2(new_n409), .A3(KEYINPUT10), .ZN(new_n410));
  INV_X1    g224(.A(new_n278), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT1), .ZN(new_n412));
  OAI22_X1  g226(.A1(new_n275), .A2(G128), .B1(new_n412), .B2(new_n265), .ZN(new_n413));
  OAI211_X1 g227(.A(new_n400), .B(new_n408), .C1(new_n411), .C2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT10), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n410), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n306), .B1(new_n405), .B2(new_n417), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n398), .A2(new_n403), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n403), .B1(new_n398), .B2(new_n400), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n307), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(new_n306), .ZN(new_n422));
  INV_X1    g236(.A(new_n417), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n385), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n414), .B1(new_n279), .B2(new_n409), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n306), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT12), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(KEYINPUT12), .A3(new_n306), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n424), .A2(new_n431), .A3(new_n385), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n382), .B(new_n189), .C1(new_n425), .C2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(KEYINPUT82), .ZN(new_n434));
  INV_X1    g248(.A(new_n385), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n405), .A2(new_n306), .A3(new_n417), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n422), .B1(new_n421), .B2(new_n423), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n424), .A2(new_n431), .A3(new_n385), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT82), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n440), .A2(new_n441), .A3(new_n382), .A4(new_n189), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n434), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n424), .A2(new_n431), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n435), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n418), .A2(new_n424), .A3(new_n385), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n382), .B1(new_n447), .B2(new_n189), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n443), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g264(.A(KEYINPUT9), .B(G234), .Z(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G221), .B1(new_n452), .B2(G902), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n453), .B(KEYINPUT79), .Z(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G214), .B1(G237), .B2(G902), .ZN(new_n457));
  OAI21_X1  g271(.A(G210), .B1(G237), .B2(G902), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n320), .B1(new_n419), .B2(new_n420), .ZN(new_n460));
  XNOR2_X1  g274(.A(G110), .B(G122), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT83), .ZN(new_n462));
  OR3_X1    g276(.A1(new_n314), .A2(new_n462), .A3(KEYINPUT5), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n314), .A2(new_n316), .A3(KEYINPUT5), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n462), .B1(new_n314), .B2(KEYINPUT5), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n463), .A2(G113), .A3(new_n464), .A4(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n409), .A2(new_n319), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n460), .A2(new_n461), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n409), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n319), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT85), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(new_n467), .ZN(new_n472));
  INV_X1    g286(.A(new_n467), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT85), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n461), .B(KEYINPUT8), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n271), .A2(new_n276), .A3(new_n194), .A4(new_n278), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n300), .A2(G125), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(G224), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n480), .A2(G953), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n481), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n477), .A2(new_n478), .A3(KEYINPUT7), .A4(new_n483), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT7), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n479), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n468), .A2(new_n476), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n189), .ZN(new_n489));
  XNOR2_X1  g303(.A(new_n479), .B(new_n481), .ZN(new_n490));
  NAND2_X1  g304(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n402), .A2(new_n404), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n473), .B1(new_n492), .B2(new_n320), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n491), .B1(new_n493), .B2(new_n461), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n460), .A2(new_n467), .ZN(new_n495));
  INV_X1    g309(.A(new_n461), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n495), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n494), .A2(new_n468), .A3(new_n497), .ZN(new_n498));
  AOI211_X1 g312(.A(new_n459), .B(new_n489), .C1(new_n490), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n490), .ZN(new_n500));
  INV_X1    g314(.A(new_n489), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n458), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n457), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n456), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT88), .ZN(new_n505));
  AOI21_X1  g319(.A(G237), .B1(new_n220), .B2(new_n222), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n506), .A2(G143), .A3(G214), .ZN(new_n507));
  AOI21_X1  g321(.A(G143), .B1(new_n506), .B2(G214), .ZN(new_n508));
  OAI21_X1  g322(.A(G131), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT17), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n223), .A2(G214), .A3(new_n322), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(new_n264), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n506), .A2(G143), .A3(G214), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n280), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n509), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n203), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n280), .B1(new_n512), .B2(new_n513), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(KEYINPUT17), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  XOR2_X1   g333(.A(G113), .B(G122), .Z(new_n520));
  XNOR2_X1  g334(.A(new_n520), .B(KEYINPUT87), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(new_n406), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n523));
  OAI211_X1 g337(.A(new_n512), .B(new_n513), .C1(new_n523), .C2(new_n280), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n240), .A2(new_n199), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n195), .A2(new_n197), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n525), .B1(new_n199), .B2(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n524), .B(new_n527), .C1(new_n509), .C2(new_n523), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n519), .A2(new_n522), .A3(new_n528), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n240), .A2(KEYINPUT19), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT19), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n531), .B1(new_n195), .B2(new_n197), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(G146), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(KEYINPUT86), .B1(new_n534), .B2(new_n239), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n240), .A2(KEYINPUT19), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n199), .B1(new_n536), .B2(new_n532), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT86), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n201), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n514), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n535), .B(new_n539), .C1(new_n517), .C2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n522), .B1(new_n541), .B2(new_n528), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n505), .B1(new_n529), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n539), .B1(new_n540), .B2(new_n517), .ZN(new_n544));
  INV_X1    g358(.A(new_n535), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n528), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n522), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n519), .A2(new_n522), .A3(new_n528), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(KEYINPUT88), .A3(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(G475), .A2(G902), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n543), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT20), .ZN(new_n553));
  NOR3_X1   g367(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n554), .B1(new_n529), .B2(new_n542), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n557), .A2(G128), .A3(new_n264), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n264), .A2(G128), .ZN(new_n559));
  INV_X1    g373(.A(G128), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G143), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n558), .B(G134), .C1(new_n562), .C2(new_n557), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT90), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(new_n559), .B2(new_n561), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n559), .A2(new_n561), .A3(new_n564), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(new_n567), .A3(new_n294), .ZN(new_n568));
  XNOR2_X1  g382(.A(G116), .B(G122), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(new_n387), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n563), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n567), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n290), .B1(new_n573), .B2(new_n565), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(G122), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(G116), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n387), .B1(new_n577), .B2(KEYINPUT14), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(new_n569), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(KEYINPUT91), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT91), .B1(new_n575), .B2(new_n579), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n572), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n451), .A2(G217), .A3(new_n219), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n294), .B1(new_n566), .B2(new_n567), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n573), .A2(new_n290), .A3(new_n565), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n579), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT91), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n580), .ZN(new_n591));
  INV_X1    g405(.A(new_n584), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n572), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(G902), .B1(new_n585), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G478), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(KEYINPUT15), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n594), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n519), .A2(new_n528), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(new_n547), .ZN(new_n599));
  AOI21_X1  g413(.A(G902), .B1(new_n599), .B2(new_n549), .ZN(new_n600));
  INV_X1    g414(.A(G475), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n223), .ZN(new_n604));
  NAND2_X1  g418(.A1(G234), .A2(G237), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n604), .A2(G902), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT21), .B(G898), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT92), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AND3_X1   g423(.A1(new_n605), .A2(G952), .A3(new_n219), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n556), .A2(new_n597), .A3(new_n603), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(KEYINPUT93), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n602), .B1(new_n553), .B2(new_n555), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT93), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n615), .A2(new_n616), .A3(new_n597), .A4(new_n612), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n381), .A2(new_n504), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G101), .ZN(G3));
  INV_X1    g434(.A(G472), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n347), .B2(new_n189), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n349), .ZN(new_n624));
  NOR3_X1   g438(.A1(new_n456), .A2(new_n261), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n500), .A2(new_n501), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n459), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n500), .A2(new_n458), .A3(new_n501), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(KEYINPUT94), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT33), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n592), .B1(new_n591), .B2(new_n572), .ZN(new_n631));
  AOI211_X1 g445(.A(new_n571), .B(new_n584), .C1(new_n590), .C2(new_n580), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n585), .A2(KEYINPUT33), .A3(new_n593), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT95), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n635), .A2(new_n636), .A3(G478), .A4(new_n189), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n633), .A2(new_n634), .A3(G478), .A4(new_n189), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT95), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT96), .B(G478), .Z(new_n641));
  OR3_X1    g455(.A1(new_n594), .A2(KEYINPUT97), .A3(new_n641), .ZN(new_n642));
  OAI21_X1  g456(.A(KEYINPUT97), .B1(new_n594), .B2(new_n641), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n615), .B1(new_n640), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT94), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n500), .A2(new_n646), .A3(new_n458), .A4(new_n501), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n647), .A2(new_n457), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n629), .A2(new_n645), .A3(new_n648), .A4(new_n612), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT98), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n625), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(new_n653), .B(KEYINPUT99), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT34), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(new_n406), .ZN(G6));
  XNOR2_X1  g470(.A(new_n602), .B(KEYINPUT100), .ZN(new_n657));
  INV_X1    g471(.A(new_n597), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n543), .A2(new_n550), .ZN(new_n659));
  INV_X1    g473(.A(new_n554), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n553), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AND3_X1   g475(.A1(new_n657), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n662), .A2(new_n629), .A3(new_n648), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n612), .B(KEYINPUT101), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n625), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT35), .B(G107), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G9));
  NOR3_X1   g482(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT36), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n669), .A2(new_n247), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n247), .ZN(new_n671));
  AND4_X1   g485(.A1(new_n189), .A2(new_n670), .A3(new_n191), .A4(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n672), .A2(new_n254), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n624), .A2(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n448), .B1(new_n434), .B2(new_n442), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n675), .A2(new_n454), .ZN(new_n676));
  INV_X1    g490(.A(new_n503), .ZN(new_n677));
  AND4_X1   g491(.A1(new_n618), .A2(new_n674), .A3(new_n676), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT37), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G110), .ZN(G12));
  INV_X1    g494(.A(KEYINPUT103), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n349), .A2(KEYINPUT32), .ZN(new_n682));
  AOI22_X1  g496(.A1(new_n682), .A2(new_n352), .B1(KEYINPUT69), .B2(new_n349), .ZN(new_n683));
  INV_X1    g497(.A(new_n356), .ZN(new_n684));
  AND3_X1   g498(.A1(new_n371), .A2(new_n358), .A3(new_n189), .ZN(new_n685));
  INV_X1    g499(.A(new_n377), .ZN(new_n686));
  NOR3_X1   g500(.A1(new_n685), .A2(new_n372), .A3(new_n686), .ZN(new_n687));
  OAI22_X1  g501(.A1(new_n683), .A2(new_n684), .B1(new_n687), .B2(new_n621), .ZN(new_n688));
  INV_X1    g502(.A(new_n673), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n647), .A2(new_n457), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n499), .A2(new_n502), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n691), .B1(new_n692), .B2(KEYINPUT94), .ZN(new_n693));
  INV_X1    g507(.A(G900), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n606), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g509(.A1(new_n695), .A2(KEYINPUT102), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(KEYINPUT102), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n696), .A2(new_n611), .A3(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n675), .A2(new_n454), .A3(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n693), .A2(new_n700), .A3(new_n662), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n681), .B1(new_n690), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n673), .B1(new_n357), .B2(new_n380), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n703), .A2(new_n663), .A3(KEYINPUT103), .A4(new_n700), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G128), .ZN(G30));
  NOR2_X1   g520(.A1(new_n615), .A2(new_n597), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n698), .B(KEYINPUT39), .Z(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n676), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n707), .B1(new_n710), .B2(KEYINPUT40), .ZN(new_n711));
  INV_X1    g525(.A(new_n457), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n692), .B(KEYINPUT38), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(KEYINPUT40), .B2(new_n710), .ZN(new_n715));
  INV_X1    g529(.A(new_n368), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n336), .B1(new_n332), .B2(new_n716), .ZN(new_n717));
  AND2_X1   g531(.A1(new_n717), .A2(new_n189), .ZN(new_n718));
  OAI22_X1  g532(.A1(new_n683), .A2(new_n684), .B1(new_n621), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n713), .A2(new_n715), .A3(new_n673), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G143), .ZN(G45));
  AND3_X1   g535(.A1(new_n629), .A2(new_n645), .A3(new_n648), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n722), .A2(new_n688), .A3(new_n689), .A4(new_n700), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G146), .ZN(G48));
  NAND2_X1  g538(.A1(new_n440), .A2(new_n189), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(G469), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n443), .A2(new_n455), .A3(new_n726), .ZN(new_n727));
  AOI211_X1 g541(.A(new_n727), .B(new_n261), .C1(new_n357), .C2(new_n380), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n728), .B1(new_n651), .B2(new_n652), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT104), .ZN(new_n730));
  XNOR2_X1  g544(.A(KEYINPUT41), .B(G113), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(G15));
  INV_X1    g546(.A(new_n727), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n381), .A2(new_n663), .A3(new_n665), .A4(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(KEYINPUT105), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n315), .ZN(G18));
  NAND4_X1  g550(.A1(new_n703), .A2(new_n618), .A3(new_n693), .A4(new_n733), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  NAND3_X1  g552(.A1(new_n629), .A2(new_n648), .A3(new_n707), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n337), .A2(new_n346), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n362), .B(KEYINPUT106), .C1(new_n369), .C2(new_n370), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n343), .ZN(new_n742));
  NOR3_X1   g556(.A1(new_n297), .A2(new_n304), .A3(new_n366), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n334), .B1(new_n308), .B2(new_n309), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT28), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(KEYINPUT70), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n368), .A2(new_n365), .A3(KEYINPUT28), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(KEYINPUT106), .B1(new_n748), .B2(new_n362), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n740), .B1(new_n742), .B2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n348), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n254), .A2(new_n257), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n751), .A2(new_n752), .A3(new_n623), .A4(new_n665), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n739), .A2(new_n753), .A3(new_n727), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n576), .ZN(G24));
  AOI211_X1 g569(.A(new_n622), .B(new_n673), .C1(new_n750), .C2(new_n348), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n637), .A2(new_n639), .B1(new_n643), .B2(new_n642), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n757), .A2(new_n615), .A3(new_n699), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n756), .A2(new_n693), .A3(new_n733), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G125), .ZN(G27));
  NAND2_X1  g574(.A1(new_n692), .A2(new_n457), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n456), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n381), .A2(new_n762), .A3(new_n758), .ZN(new_n763));
  XNOR2_X1  g577(.A(KEYINPUT107), .B(KEYINPUT42), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n752), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n682), .A2(new_n352), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n766), .B1(new_n380), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n762), .A2(new_n768), .A3(KEYINPUT42), .A4(new_n758), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n765), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT108), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n765), .A2(KEYINPUT108), .A3(new_n769), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(KEYINPUT109), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(new_n280), .ZN(G33));
  NAND4_X1  g590(.A1(new_n381), .A2(new_n762), .A3(new_n662), .A4(new_n698), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  NAND2_X1  g592(.A1(new_n640), .A2(new_n644), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n615), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT110), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT111), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT43), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT111), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n783), .B1(new_n780), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n782), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n781), .A2(KEYINPUT111), .A3(new_n783), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n624), .A3(new_n689), .A4(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT44), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n447), .B(KEYINPUT45), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(G469), .ZN(new_n792));
  NAND2_X1  g606(.A1(G469), .A2(G902), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(KEYINPUT46), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT46), .ZN(new_n795));
  OAI211_X1 g609(.A(new_n795), .B(G469), .C1(new_n791), .C2(G902), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n794), .A2(new_n443), .A3(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n455), .A3(new_n709), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n790), .A2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n761), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n788), .B2(new_n789), .ZN(new_n802));
  OR2_X1    g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G137), .ZN(G39));
  NAND2_X1  g618(.A1(new_n797), .A2(new_n455), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT47), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n688), .A2(new_n761), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n261), .A3(new_n758), .A4(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n809), .B(G140), .ZN(G42));
  AND3_X1   g624(.A1(new_n751), .A2(new_n752), .A3(new_n623), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n786), .A2(new_n610), .A3(new_n811), .A4(new_n787), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n727), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n813), .A2(new_n712), .A3(new_n714), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n813), .A2(KEYINPUT50), .A3(new_n712), .A4(new_n714), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n812), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n443), .A2(new_n726), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n820), .A2(new_n455), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n819), .B(new_n801), .C1(new_n807), .C2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n786), .A2(new_n787), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n761), .A2(new_n727), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n823), .A2(new_n610), .A3(new_n756), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n719), .A2(new_n611), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n761), .A2(new_n261), .A3(new_n727), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n827), .A3(new_n615), .A4(new_n757), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(KEYINPUT115), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n822), .A2(new_n825), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n818), .B(new_n830), .C1(new_n831), .C2(KEYINPUT51), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n826), .A2(new_n645), .A3(new_n827), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(G952), .A3(new_n219), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n823), .A2(new_n610), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n768), .A3(new_n824), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT48), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT48), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n835), .A2(new_n838), .A3(new_n768), .A4(new_n824), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n834), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n822), .A2(new_n825), .A3(new_n829), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n816), .B2(new_n817), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT51), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n844), .B1(new_n842), .B2(KEYINPUT114), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n678), .A2(new_n754), .ZN(new_n848));
  INV_X1    g662(.A(new_n645), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n615), .A2(new_n658), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n503), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n625), .A2(new_n665), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n729), .A2(new_n848), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n737), .A2(new_n734), .A3(new_n619), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n657), .A2(new_n661), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n658), .A2(new_n699), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n703), .A2(new_n762), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n762), .A2(new_n758), .A3(new_n756), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n777), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n853), .A2(new_n854), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n723), .A2(new_n759), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(new_n702), .B2(new_n704), .ZN(new_n862));
  INV_X1    g676(.A(new_n739), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n863), .A2(new_n719), .A3(new_n673), .A4(new_n700), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT52), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n723), .A2(new_n759), .ZN(new_n866));
  AND4_X1   g680(.A1(KEYINPUT52), .A2(new_n705), .A3(new_n866), .A4(new_n864), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n774), .B(new_n860), .C1(new_n865), .C2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n765), .A2(KEYINPUT108), .A3(new_n769), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT108), .B1(new_n765), .B2(new_n769), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n859), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n737), .A2(new_n734), .A3(new_n619), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n504), .A2(new_n618), .A3(new_n674), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n863), .A2(new_n811), .A3(new_n665), .A4(new_n733), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n852), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n874), .A2(new_n875), .A3(new_n878), .A4(new_n729), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n873), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n705), .A2(new_n866), .A3(new_n864), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT52), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n705), .A2(new_n866), .A3(KEYINPUT52), .A4(new_n864), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n880), .A2(KEYINPUT53), .A3(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n870), .A2(new_n886), .A3(KEYINPUT113), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT113), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n868), .A2(new_n888), .A3(new_n869), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n887), .A2(KEYINPUT54), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n813), .A2(new_n693), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT54), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n770), .A2(KEYINPUT53), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n883), .B2(new_n884), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n894), .A2(new_n860), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n870), .A2(new_n892), .A3(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n847), .A2(new_n890), .A3(new_n891), .A4(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(G952), .B2(G953), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n820), .A2(KEYINPUT49), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n899), .B(KEYINPUT112), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n820), .A2(KEYINPUT49), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n766), .A2(new_n454), .A3(new_n712), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n714), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  OR4_X1    g717(.A1(new_n719), .A2(new_n900), .A3(new_n903), .A4(new_n780), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n898), .A2(new_n904), .ZN(G75));
  XOR2_X1   g719(.A(new_n498), .B(new_n490), .Z(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT116), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n907), .B(KEYINPUT55), .ZN(new_n908));
  AOI21_X1  g722(.A(KEYINPUT53), .B1(new_n880), .B2(new_n885), .ZN(new_n909));
  INV_X1    g723(.A(new_n893), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n885), .A2(new_n860), .A3(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(G210), .B(G902), .C1(new_n909), .C2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT56), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n908), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n223), .A2(G952), .ZN(new_n915));
  XNOR2_X1  g729(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n912), .A2(new_n908), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n917), .A2(KEYINPUT118), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT118), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n912), .A2(new_n919), .A3(new_n908), .A4(new_n916), .ZN(new_n920));
  AOI211_X1 g734(.A(new_n914), .B(new_n915), .C1(new_n918), .C2(new_n920), .ZN(G51));
  OAI21_X1  g735(.A(KEYINPUT54), .B1(new_n909), .B2(new_n911), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n923), .A3(new_n896), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n868), .A2(new_n869), .B1(new_n894), .B2(new_n860), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(KEYINPUT119), .A3(new_n892), .ZN(new_n926));
  XOR2_X1   g740(.A(new_n793), .B(KEYINPUT57), .Z(new_n927));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n440), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n925), .A2(new_n189), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n930), .A2(G469), .A3(new_n791), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n915), .B1(new_n929), .B2(new_n931), .ZN(G54));
  NAND3_X1  g746(.A1(new_n930), .A2(KEYINPUT58), .A3(G475), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n933), .A2(new_n659), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n933), .A2(new_n659), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n934), .A2(new_n935), .A3(new_n915), .ZN(G60));
  XOR2_X1   g750(.A(new_n635), .B(KEYINPUT120), .Z(new_n937));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT59), .Z(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n924), .A2(new_n926), .A3(new_n937), .A4(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n915), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n939), .B1(new_n890), .B2(new_n896), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n941), .B(new_n942), .C1(new_n943), .C2(new_n937), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(G63));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT60), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n256), .B1(new_n925), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n870), .B2(new_n895), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n670), .A2(new_n671), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT121), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT121), .ZN(new_n953));
  NOR4_X1   g767(.A1(new_n925), .A2(new_n953), .A3(new_n950), .A4(new_n947), .ZN(new_n954));
  OAI211_X1 g768(.A(new_n942), .B(new_n948), .C1(new_n952), .C2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT61), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g771(.A(new_n947), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n909), .B2(new_n911), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n953), .B1(new_n959), .B2(new_n950), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n949), .A2(KEYINPUT121), .A3(new_n951), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n962), .A2(KEYINPUT61), .A3(new_n942), .A4(new_n948), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n957), .A2(new_n963), .ZN(G66));
  OAI21_X1  g778(.A(G953), .B1(new_n608), .B2(new_n480), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n853), .A2(new_n854), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n965), .B1(new_n966), .B2(new_n604), .ZN(new_n967));
  INV_X1    g781(.A(new_n498), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n968), .B1(G898), .B2(new_n223), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT122), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n967), .B(new_n970), .ZN(G69));
  NAND2_X1  g785(.A1(new_n705), .A2(new_n866), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n972), .A2(KEYINPUT123), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT123), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n862), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n973), .A2(new_n975), .A3(new_n720), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT62), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n305), .A2(new_n310), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n530), .A2(new_n533), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n979), .B(new_n980), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n803), .A2(new_n809), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n710), .A2(new_n761), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n849), .A2(new_n850), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n983), .A2(new_n381), .A3(new_n984), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n978), .A2(new_n981), .A3(new_n982), .A4(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n799), .A2(new_n863), .A3(new_n768), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n809), .B(new_n987), .C1(new_n800), .C2(new_n802), .ZN(new_n988));
  INV_X1    g802(.A(new_n777), .ZN(new_n989));
  NOR2_X1   g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n990), .A2(new_n774), .A3(new_n973), .A4(new_n975), .ZN(new_n991));
  INV_X1    g805(.A(new_n981), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n986), .A2(new_n993), .A3(new_n223), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n992), .A2(G227), .A3(new_n604), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(KEYINPUT124), .ZN(new_n997));
  AOI21_X1  g811(.A(G227), .B1(new_n992), .B2(KEYINPUT124), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n604), .B1(new_n998), .B2(new_n694), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n999), .ZN(G72));
  NAND2_X1  g814(.A1(G472), .A2(G902), .ZN(new_n1001));
  XOR2_X1   g815(.A(new_n1001), .B(KEYINPUT63), .Z(new_n1002));
  INV_X1    g816(.A(new_n966), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1002), .B1(new_n991), .B2(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n375), .B(KEYINPUT125), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n343), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1006), .B(KEYINPUT126), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n376), .A2(new_n336), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n887), .A2(new_n889), .A3(new_n1002), .A4(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1008), .A2(new_n942), .A3(new_n1010), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n978), .A2(new_n966), .A3(new_n982), .A4(new_n985), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1005), .B1(new_n1012), .B2(new_n1002), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1011), .B1(new_n332), .B2(new_n1013), .ZN(G57));
endmodule


