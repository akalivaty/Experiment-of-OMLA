

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579;

  INV_X1 U322 ( .A(n536), .ZN(n539) );
  NOR2_X1 U323 ( .A1(n555), .A2(n498), .ZN(n499) );
  INV_X1 U324 ( .A(n537), .ZN(n538) );
  NAND2_X1 U325 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U326 ( .A(n322), .B(n321), .ZN(n328) );
  XNOR2_X1 U327 ( .A(n328), .B(n327), .ZN(n334) );
  NOR2_X1 U328 ( .A1(n546), .A2(n545), .ZN(n560) );
  XOR2_X1 U329 ( .A(n569), .B(KEYINPUT41), .Z(n552) );
  XOR2_X1 U330 ( .A(n543), .B(KEYINPUT28), .Z(n514) );
  XNOR2_X1 U331 ( .A(KEYINPUT2), .B(KEYINPUT87), .ZN(n290) );
  XNOR2_X1 U332 ( .A(n290), .B(KEYINPUT3), .ZN(n291) );
  XOR2_X1 U333 ( .A(n291), .B(KEYINPUT86), .Z(n293) );
  XNOR2_X1 U334 ( .A(G141GAT), .B(G155GAT), .ZN(n292) );
  XNOR2_X1 U335 ( .A(n293), .B(n292), .ZN(n398) );
  XOR2_X1 U336 ( .A(G57GAT), .B(G148GAT), .Z(n295) );
  XNOR2_X1 U337 ( .A(G1GAT), .B(G127GAT), .ZN(n294) );
  XNOR2_X1 U338 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U339 ( .A(KEYINPUT92), .B(KEYINPUT93), .Z(n297) );
  XNOR2_X1 U340 ( .A(KEYINPUT95), .B(KEYINPUT94), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U342 ( .A(n299), .B(n298), .Z(n306) );
  XOR2_X1 U343 ( .A(G120GAT), .B(KEYINPUT0), .Z(n301) );
  XNOR2_X1 U344 ( .A(G113GAT), .B(KEYINPUT78), .ZN(n300) );
  XNOR2_X1 U345 ( .A(n301), .B(n300), .ZN(n358) );
  XOR2_X1 U346 ( .A(G85GAT), .B(G162GAT), .Z(n303) );
  XNOR2_X1 U347 ( .A(G29GAT), .B(G134GAT), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U349 ( .A(n358), .B(n304), .ZN(n305) );
  XNOR2_X1 U350 ( .A(n306), .B(n305), .ZN(n313) );
  XOR2_X1 U351 ( .A(KEYINPUT91), .B(KEYINPUT4), .Z(n308) );
  XNOR2_X1 U352 ( .A(KEYINPUT96), .B(KEYINPUT97), .ZN(n307) );
  XNOR2_X1 U353 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U354 ( .A(KEYINPUT5), .B(n309), .Z(n311) );
  NAND2_X1 U355 ( .A1(G225GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U356 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U357 ( .A(n313), .B(n312), .Z(n315) );
  XNOR2_X1 U358 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n314) );
  XNOR2_X1 U359 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U360 ( .A(n398), .B(n316), .ZN(n542) );
  XOR2_X1 U361 ( .A(KEYINPUT74), .B(KEYINPUT73), .Z(n318) );
  NAND2_X1 U362 ( .A1(G230GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U363 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U364 ( .A(KEYINPUT33), .B(n319), .ZN(n322) );
  XNOR2_X1 U365 ( .A(G99GAT), .B(G85GAT), .ZN(n320) );
  XNOR2_X1 U366 ( .A(n320), .B(KEYINPUT72), .ZN(n416) );
  INV_X1 U367 ( .A(n416), .ZN(n321) );
  XOR2_X1 U368 ( .A(KEYINPUT71), .B(KEYINPUT32), .Z(n324) );
  XNOR2_X1 U369 ( .A(G120GAT), .B(KEYINPUT31), .ZN(n323) );
  XNOR2_X1 U370 ( .A(n324), .B(n323), .ZN(n326) );
  XNOR2_X1 U371 ( .A(G176GAT), .B(G92GAT), .ZN(n325) );
  XNOR2_X1 U372 ( .A(n325), .B(G64GAT), .ZN(n378) );
  XOR2_X1 U373 ( .A(n326), .B(n378), .Z(n327) );
  XNOR2_X1 U374 ( .A(G106GAT), .B(G204GAT), .ZN(n329) );
  XNOR2_X1 U375 ( .A(n329), .B(G148GAT), .ZN(n390) );
  XOR2_X1 U376 ( .A(KEYINPUT13), .B(KEYINPUT70), .Z(n331) );
  XNOR2_X1 U377 ( .A(G71GAT), .B(G78GAT), .ZN(n330) );
  XNOR2_X1 U378 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U379 ( .A(G57GAT), .B(n332), .Z(n440) );
  XNOR2_X1 U380 ( .A(n390), .B(n440), .ZN(n333) );
  XNOR2_X1 U381 ( .A(n334), .B(n333), .ZN(n569) );
  XOR2_X1 U382 ( .A(G1GAT), .B(G8GAT), .Z(n336) );
  XNOR2_X1 U383 ( .A(G22GAT), .B(G15GAT), .ZN(n335) );
  XNOR2_X1 U384 ( .A(n336), .B(n335), .ZN(n429) );
  XOR2_X1 U385 ( .A(n429), .B(KEYINPUT68), .Z(n338) );
  NAND2_X1 U386 ( .A1(G229GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U387 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U388 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n340) );
  XNOR2_X1 U389 ( .A(KEYINPUT29), .B(KEYINPUT30), .ZN(n339) );
  XNOR2_X1 U390 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U391 ( .A(n342), .B(n341), .Z(n351) );
  XNOR2_X1 U392 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n343) );
  XNOR2_X1 U393 ( .A(n343), .B(G29GAT), .ZN(n344) );
  XOR2_X1 U394 ( .A(n344), .B(KEYINPUT8), .Z(n346) );
  XNOR2_X1 U395 ( .A(G43GAT), .B(G50GAT), .ZN(n345) );
  XNOR2_X1 U396 ( .A(n346), .B(n345), .ZN(n426) );
  XOR2_X1 U397 ( .A(G113GAT), .B(G141GAT), .Z(n348) );
  XNOR2_X1 U398 ( .A(G169GAT), .B(G197GAT), .ZN(n347) );
  XNOR2_X1 U399 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U400 ( .A(n426), .B(n349), .ZN(n350) );
  XNOR2_X1 U401 ( .A(n351), .B(n350), .ZN(n565) );
  XOR2_X1 U402 ( .A(n565), .B(KEYINPUT69), .Z(n547) );
  INV_X1 U403 ( .A(n547), .ZN(n504) );
  NOR2_X1 U404 ( .A1(n569), .A2(n504), .ZN(n460) );
  XOR2_X1 U405 ( .A(KEYINPUT101), .B(KEYINPUT25), .Z(n403) );
  XOR2_X1 U406 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n353) );
  XNOR2_X1 U407 ( .A(G71GAT), .B(KEYINPUT79), .ZN(n352) );
  XNOR2_X1 U408 ( .A(n353), .B(n352), .ZN(n368) );
  XOR2_X1 U409 ( .A(G183GAT), .B(G127GAT), .Z(n430) );
  XOR2_X1 U410 ( .A(G99GAT), .B(n430), .Z(n355) );
  XOR2_X1 U411 ( .A(G190GAT), .B(G134GAT), .Z(n419) );
  XNOR2_X1 U412 ( .A(G43GAT), .B(n419), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n364) );
  XOR2_X1 U414 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n357) );
  XNOR2_X1 U415 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n356) );
  XNOR2_X1 U416 ( .A(n357), .B(n356), .ZN(n379) );
  XNOR2_X1 U417 ( .A(n358), .B(n379), .ZN(n362) );
  XOR2_X1 U418 ( .A(G176GAT), .B(KEYINPUT80), .Z(n360) );
  XNOR2_X1 U419 ( .A(G15GAT), .B(KEYINPUT20), .ZN(n359) );
  XNOR2_X1 U420 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U421 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U422 ( .A(n364), .B(n363), .Z(n366) );
  NAND2_X1 U423 ( .A1(G227GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U425 ( .A(n368), .B(n367), .ZN(n546) );
  XOR2_X1 U426 ( .A(KEYINPUT21), .B(KEYINPUT85), .Z(n370) );
  XNOR2_X1 U427 ( .A(KEYINPUT84), .B(G211GAT), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U429 ( .A(G197GAT), .B(n371), .Z(n393) );
  XOR2_X1 U430 ( .A(G204GAT), .B(G183GAT), .Z(n373) );
  XNOR2_X1 U431 ( .A(G8GAT), .B(G190GAT), .ZN(n372) );
  XNOR2_X1 U432 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U433 ( .A(G218GAT), .B(G36GAT), .Z(n375) );
  NAND2_X1 U434 ( .A1(G226GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U436 ( .A(n377), .B(n376), .Z(n381) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n393), .B(n382), .ZN(n537) );
  NOR2_X1 U440 ( .A1(n546), .A2(n537), .ZN(n383) );
  XOR2_X1 U441 ( .A(KEYINPUT100), .B(n383), .Z(n401) );
  XOR2_X1 U442 ( .A(G218GAT), .B(G162GAT), .Z(n418) );
  XOR2_X1 U443 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n385) );
  XNOR2_X1 U444 ( .A(G50GAT), .B(G78GAT), .ZN(n384) );
  XNOR2_X1 U445 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U446 ( .A(n418), .B(n386), .Z(n388) );
  NAND2_X1 U447 ( .A1(G228GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U449 ( .A(n389), .B(KEYINPUT83), .Z(n392) );
  XNOR2_X1 U450 ( .A(n390), .B(KEYINPUT90), .ZN(n391) );
  XNOR2_X1 U451 ( .A(n392), .B(n391), .ZN(n397) );
  XOR2_X1 U452 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n395) );
  XNOR2_X1 U453 ( .A(n393), .B(KEYINPUT88), .ZN(n394) );
  XNOR2_X1 U454 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U455 ( .A(n397), .B(n396), .Z(n400) );
  XNOR2_X1 U456 ( .A(G22GAT), .B(n398), .ZN(n399) );
  XNOR2_X1 U457 ( .A(n400), .B(n399), .ZN(n543) );
  NAND2_X1 U458 ( .A1(n401), .A2(n543), .ZN(n402) );
  XNOR2_X1 U459 ( .A(n403), .B(n402), .ZN(n407) );
  INV_X1 U460 ( .A(n546), .ZN(n487) );
  NOR2_X1 U461 ( .A1(n487), .A2(n543), .ZN(n404) );
  XNOR2_X1 U462 ( .A(KEYINPUT26), .B(n404), .ZN(n564) );
  XNOR2_X1 U463 ( .A(KEYINPUT27), .B(KEYINPUT98), .ZN(n405) );
  XOR2_X1 U464 ( .A(n405), .B(n537), .Z(n409) );
  AND2_X1 U465 ( .A1(n564), .A2(n409), .ZN(n406) );
  NOR2_X1 U466 ( .A1(n407), .A2(n406), .ZN(n408) );
  NOR2_X1 U467 ( .A1(n408), .A2(n542), .ZN(n413) );
  NAND2_X1 U468 ( .A1(n542), .A2(n409), .ZN(n410) );
  XOR2_X1 U469 ( .A(n410), .B(KEYINPUT99), .Z(n511) );
  OR2_X1 U470 ( .A1(n487), .A2(n511), .ZN(n411) );
  NOR2_X1 U471 ( .A1(n514), .A2(n411), .ZN(n412) );
  NOR2_X1 U472 ( .A1(n413), .A2(n412), .ZN(n456) );
  XOR2_X1 U473 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n415) );
  XNOR2_X1 U474 ( .A(KEYINPUT9), .B(KEYINPUT75), .ZN(n414) );
  XNOR2_X1 U475 ( .A(n415), .B(n414), .ZN(n417) );
  XOR2_X1 U476 ( .A(n417), .B(n416), .Z(n421) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U479 ( .A(G92GAT), .B(KEYINPUT65), .Z(n423) );
  NAND2_X1 U480 ( .A1(G232GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U481 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U482 ( .A(n425), .B(n424), .Z(n428) );
  XNOR2_X1 U483 ( .A(n426), .B(G106GAT), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n496) );
  INV_X1 U485 ( .A(n496), .ZN(n559) );
  XOR2_X1 U486 ( .A(n430), .B(n429), .Z(n432) );
  NAND2_X1 U487 ( .A1(G231GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U489 ( .A(KEYINPUT76), .B(KEYINPUT15), .Z(n434) );
  XNOR2_X1 U490 ( .A(KEYINPUT77), .B(KEYINPUT12), .ZN(n433) );
  XNOR2_X1 U491 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U492 ( .A(n436), .B(n435), .Z(n442) );
  XOR2_X1 U493 ( .A(KEYINPUT14), .B(G64GAT), .Z(n438) );
  XNOR2_X1 U494 ( .A(G155GAT), .B(G211GAT), .ZN(n437) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n573) );
  INV_X1 U498 ( .A(n573), .ZN(n500) );
  NOR2_X1 U499 ( .A1(n559), .A2(n500), .ZN(n443) );
  XOR2_X1 U500 ( .A(KEYINPUT16), .B(n443), .Z(n444) );
  NOR2_X1 U501 ( .A1(n456), .A2(n444), .ZN(n470) );
  AND2_X1 U502 ( .A1(n460), .A2(n470), .ZN(n451) );
  NAND2_X1 U503 ( .A1(n542), .A2(n451), .ZN(n445) );
  XNOR2_X1 U504 ( .A(n445), .B(KEYINPUT34), .ZN(n446) );
  XNOR2_X1 U505 ( .A(G1GAT), .B(n446), .ZN(G1324GAT) );
  NAND2_X1 U506 ( .A1(n451), .A2(n538), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n447), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U508 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n449) );
  NAND2_X1 U509 ( .A1(n451), .A2(n487), .ZN(n448) );
  XNOR2_X1 U510 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U511 ( .A(G15GAT), .B(n450), .ZN(G1326GAT) );
  NAND2_X1 U512 ( .A1(n451), .A2(n514), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n452), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U514 ( .A(KEYINPUT103), .B(KEYINPUT39), .Z(n454) );
  XNOR2_X1 U515 ( .A(G29GAT), .B(KEYINPUT106), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n454), .B(n453), .ZN(n463) );
  XNOR2_X1 U517 ( .A(n496), .B(KEYINPUT104), .ZN(n455) );
  XNOR2_X1 U518 ( .A(n455), .B(KEYINPUT36), .ZN(n577) );
  NOR2_X1 U519 ( .A1(n573), .A2(n456), .ZN(n457) );
  XNOR2_X1 U520 ( .A(n457), .B(KEYINPUT105), .ZN(n458) );
  NOR2_X1 U521 ( .A1(n577), .A2(n458), .ZN(n459) );
  XOR2_X1 U522 ( .A(KEYINPUT37), .B(n459), .Z(n481) );
  NAND2_X1 U523 ( .A1(n481), .A2(n460), .ZN(n461) );
  XOR2_X1 U524 ( .A(KEYINPUT38), .B(n461), .Z(n467) );
  NAND2_X1 U525 ( .A1(n467), .A2(n542), .ZN(n462) );
  XOR2_X1 U526 ( .A(n463), .B(n462), .Z(G1328GAT) );
  NAND2_X1 U527 ( .A1(n538), .A2(n467), .ZN(n464) );
  XNOR2_X1 U528 ( .A(G36GAT), .B(n464), .ZN(G1329GAT) );
  NAND2_X1 U529 ( .A1(n467), .A2(n487), .ZN(n465) );
  XNOR2_X1 U530 ( .A(n465), .B(KEYINPUT40), .ZN(n466) );
  XNOR2_X1 U531 ( .A(G43GAT), .B(n466), .ZN(G1330GAT) );
  NAND2_X1 U532 ( .A1(n467), .A2(n514), .ZN(n468) );
  XNOR2_X1 U533 ( .A(n468), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT42), .B(KEYINPUT107), .Z(n472) );
  INV_X1 U535 ( .A(n552), .ZN(n469) );
  NOR2_X1 U536 ( .A1(n565), .A2(n469), .ZN(n482) );
  AND2_X1 U537 ( .A1(n482), .A2(n470), .ZN(n477) );
  NAND2_X1 U538 ( .A1(n477), .A2(n542), .ZN(n471) );
  XNOR2_X1 U539 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U540 ( .A(G57GAT), .B(n473), .ZN(G1332GAT) );
  NAND2_X1 U541 ( .A1(n477), .A2(n538), .ZN(n474) );
  XNOR2_X1 U542 ( .A(n474), .B(KEYINPUT108), .ZN(n475) );
  XNOR2_X1 U543 ( .A(G64GAT), .B(n475), .ZN(G1333GAT) );
  NAND2_X1 U544 ( .A1(n477), .A2(n487), .ZN(n476) );
  XNOR2_X1 U545 ( .A(n476), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n479) );
  NAND2_X1 U547 ( .A1(n477), .A2(n514), .ZN(n478) );
  XNOR2_X1 U548 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U549 ( .A(G78GAT), .B(n480), .Z(G1335GAT) );
  XOR2_X1 U550 ( .A(G85GAT), .B(KEYINPUT111), .Z(n485) );
  NAND2_X1 U551 ( .A1(n482), .A2(n481), .ZN(n483) );
  XOR2_X1 U552 ( .A(KEYINPUT110), .B(n483), .Z(n491) );
  NAND2_X1 U553 ( .A1(n491), .A2(n542), .ZN(n484) );
  XNOR2_X1 U554 ( .A(n485), .B(n484), .ZN(G1336GAT) );
  NAND2_X1 U555 ( .A1(n491), .A2(n538), .ZN(n486) );
  XNOR2_X1 U556 ( .A(n486), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n489) );
  NAND2_X1 U558 ( .A1(n487), .A2(n491), .ZN(n488) );
  XNOR2_X1 U559 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U560 ( .A(G99GAT), .B(n490), .ZN(G1338GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT44), .B(KEYINPUT114), .Z(n493) );
  NAND2_X1 U562 ( .A1(n514), .A2(n491), .ZN(n492) );
  XNOR2_X1 U563 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U564 ( .A(G106GAT), .B(n494), .Z(G1339GAT) );
  XNOR2_X1 U565 ( .A(KEYINPUT64), .B(KEYINPUT117), .ZN(n510) );
  XOR2_X1 U566 ( .A(n573), .B(KEYINPUT115), .Z(n555) );
  NAND2_X1 U567 ( .A1(n565), .A2(n552), .ZN(n495) );
  XNOR2_X1 U568 ( .A(KEYINPUT46), .B(n495), .ZN(n497) );
  NAND2_X1 U569 ( .A1(n497), .A2(n496), .ZN(n498) );
  XNOR2_X1 U570 ( .A(KEYINPUT47), .B(n499), .ZN(n507) );
  NOR2_X1 U571 ( .A1(n577), .A2(n500), .ZN(n501) );
  XOR2_X1 U572 ( .A(KEYINPUT45), .B(n501), .Z(n502) );
  NOR2_X1 U573 ( .A1(n569), .A2(n502), .ZN(n503) );
  XNOR2_X1 U574 ( .A(n503), .B(KEYINPUT116), .ZN(n505) );
  NAND2_X1 U575 ( .A1(n505), .A2(n504), .ZN(n506) );
  NAND2_X1 U576 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U577 ( .A(n508), .B(KEYINPUT48), .ZN(n509) );
  XNOR2_X1 U578 ( .A(n510), .B(n509), .ZN(n536) );
  NOR2_X1 U579 ( .A1(n536), .A2(n511), .ZN(n512) );
  XOR2_X1 U580 ( .A(KEYINPUT118), .B(n512), .Z(n524) );
  OR2_X1 U581 ( .A1(n546), .A2(n524), .ZN(n513) );
  NOR2_X1 U582 ( .A1(n514), .A2(n513), .ZN(n521) );
  NAND2_X1 U583 ( .A1(n547), .A2(n521), .ZN(n515) );
  XNOR2_X1 U584 ( .A(G113GAT), .B(n515), .ZN(G1340GAT) );
  XOR2_X1 U585 ( .A(G120GAT), .B(KEYINPUT49), .Z(n517) );
  NAND2_X1 U586 ( .A1(n521), .A2(n552), .ZN(n516) );
  XNOR2_X1 U587 ( .A(n517), .B(n516), .ZN(G1341GAT) );
  XOR2_X1 U588 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n519) );
  NAND2_X1 U589 ( .A1(n521), .A2(n555), .ZN(n518) );
  XNOR2_X1 U590 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U591 ( .A(G127GAT), .B(n520), .ZN(G1342GAT) );
  XOR2_X1 U592 ( .A(G134GAT), .B(KEYINPUT51), .Z(n523) );
  NAND2_X1 U593 ( .A1(n521), .A2(n559), .ZN(n522) );
  XNOR2_X1 U594 ( .A(n523), .B(n522), .ZN(G1343GAT) );
  INV_X1 U595 ( .A(n564), .ZN(n525) );
  NOR2_X1 U596 ( .A1(n525), .A2(n524), .ZN(n533) );
  NAND2_X1 U597 ( .A1(n565), .A2(n533), .ZN(n526) );
  XNOR2_X1 U598 ( .A(KEYINPUT120), .B(n526), .ZN(n527) );
  XNOR2_X1 U599 ( .A(G141GAT), .B(n527), .ZN(G1344GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n529) );
  NAND2_X1 U601 ( .A1(n533), .A2(n552), .ZN(n528) );
  XNOR2_X1 U602 ( .A(n529), .B(n528), .ZN(n531) );
  XOR2_X1 U603 ( .A(G148GAT), .B(KEYINPUT121), .Z(n530) );
  XNOR2_X1 U604 ( .A(n531), .B(n530), .ZN(G1345GAT) );
  NAND2_X1 U605 ( .A1(n533), .A2(n573), .ZN(n532) );
  XNOR2_X1 U606 ( .A(n532), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U607 ( .A1(n559), .A2(n533), .ZN(n534) );
  XNOR2_X1 U608 ( .A(n534), .B(KEYINPUT122), .ZN(n535) );
  XNOR2_X1 U609 ( .A(G162GAT), .B(n535), .ZN(G1347GAT) );
  XNOR2_X1 U610 ( .A(n540), .B(KEYINPUT54), .ZN(n541) );
  NOR2_X1 U611 ( .A1(n542), .A2(n541), .ZN(n563) );
  NAND2_X1 U612 ( .A1(n543), .A2(n563), .ZN(n544) );
  XOR2_X1 U613 ( .A(KEYINPUT55), .B(n544), .Z(n545) );
  NAND2_X1 U614 ( .A1(n560), .A2(n547), .ZN(n548) );
  XNOR2_X1 U615 ( .A(n548), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n550) );
  XNOR2_X1 U617 ( .A(G176GAT), .B(KEYINPUT123), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(n551) );
  XOR2_X1 U619 ( .A(KEYINPUT56), .B(n551), .Z(n554) );
  NAND2_X1 U620 ( .A1(n560), .A2(n552), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(G1349GAT) );
  NAND2_X1 U622 ( .A1(n560), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U624 ( .A(G190GAT), .B(KEYINPUT126), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n557), .B(KEYINPUT125), .ZN(n558) );
  XOR2_X1 U626 ( .A(KEYINPUT58), .B(n558), .Z(n562) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(G1351GAT) );
  XOR2_X1 U629 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n567) );
  NAND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n576) );
  INV_X1 U631 ( .A(n576), .ZN(n574) );
  NAND2_X1 U632 ( .A1(n574), .A2(n565), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT61), .B(KEYINPUT127), .Z(n571) );
  NAND2_X1 U636 ( .A1(n574), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(G204GAT), .B(n572), .Z(G1353GAT) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U641 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U642 ( .A(KEYINPUT62), .B(n578), .Z(n579) );
  XNOR2_X1 U643 ( .A(G218GAT), .B(n579), .ZN(G1355GAT) );
endmodule

