//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n890, new_n891, new_n893, new_n894, new_n895, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n954, new_n955, new_n956, new_n957, new_n959, new_n960;
  INV_X1    g000(.A(G183gat), .ZN(new_n202));
  OAI21_X1  g001(.A(KEYINPUT27), .B1(new_n202), .B2(KEYINPUT65), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT65), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT27), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n204), .A2(new_n205), .A3(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT28), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT27), .B(G183gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(KEYINPUT28), .A3(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G169gat), .ZN(new_n214));
  INV_X1    g013(.A(G176gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT26), .ZN(new_n216));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n214), .A2(new_n215), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT26), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G169gat), .B2(G176gat), .ZN(new_n220));
  OAI211_X1 g019(.A(new_n216), .B(new_n217), .C1(new_n218), .C2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n213), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n217), .A2(KEYINPUT24), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n225), .A2(G183gat), .A3(G190gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n224), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n202), .A2(new_n207), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n218), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  OR3_X1    g028(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  AND3_X1   g031(.A1(new_n229), .A2(KEYINPUT25), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT25), .B1(new_n229), .B2(new_n232), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n223), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G120gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G113gat), .ZN(new_n237));
  INV_X1    g036(.A(G113gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n238), .A2(G120gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n241));
  INV_X1    g040(.A(G134gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(G127gat), .ZN(new_n243));
  INV_X1    g042(.A(G127gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G134gat), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n240), .A2(new_n241), .A3(new_n243), .A4(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n245), .ZN(new_n247));
  XNOR2_X1  g046(.A(G113gat), .B(G120gat), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n247), .B1(new_n248), .B2(KEYINPUT1), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n246), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n221), .B1(new_n210), .B2(new_n212), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n225), .B1(G183gat), .B2(G190gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n217), .A2(KEYINPUT24), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n228), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n218), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(new_n232), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT25), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n229), .A2(KEYINPUT25), .A3(new_n232), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n252), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g060(.A1(new_n246), .A2(new_n249), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G227gat), .A2(G233gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n251), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(KEYINPUT34), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT34), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n264), .B(KEYINPUT64), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n251), .A2(new_n263), .A3(new_n267), .A4(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G71gat), .B(G99gat), .ZN(new_n272));
  INV_X1    g071(.A(G43gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(KEYINPUT66), .B(G15gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n268), .B1(new_n251), .B2(new_n263), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT32), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n278), .A2(KEYINPUT33), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI211_X1 g081(.A(KEYINPUT67), .B(new_n276), .C1(new_n277), .C2(new_n279), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n276), .A2(KEYINPUT33), .ZN(new_n285));
  NOR3_X1   g084(.A1(new_n277), .A2(new_n278), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n271), .B1(new_n284), .B2(new_n287), .ZN(new_n288));
  AOI211_X1 g087(.A(new_n286), .B(new_n270), .C1(new_n282), .C2(new_n283), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT68), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT36), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(KEYINPUT68), .B(KEYINPUT36), .C1(new_n288), .C2(new_n289), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(KEYINPUT77), .B(KEYINPUT0), .Z(new_n295));
  XNOR2_X1  g094(.A(G1gat), .B(G29gat), .ZN(new_n296));
  XNOR2_X1  g095(.A(new_n295), .B(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G57gat), .B(G85gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(KEYINPUT2), .ZN(new_n301));
  INV_X1    g100(.A(G141gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(G148gat), .ZN(new_n303));
  INV_X1    g102(.A(G148gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(new_n304), .A2(G141gat), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n301), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT75), .ZN(new_n307));
  XNOR2_X1  g106(.A(new_n300), .B(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G155gat), .ZN(new_n309));
  INV_X1    g108(.A(G162gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n306), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT76), .B1(new_n303), .B2(new_n305), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n300), .B1(new_n311), .B2(KEYINPUT2), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n304), .A2(G141gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n302), .A2(G148gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT76), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n313), .A2(new_n314), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n312), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(KEYINPUT4), .B1(new_n320), .B2(new_n250), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT4), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n262), .A2(new_n322), .A3(new_n312), .A4(new_n319), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G225gat), .A2(G233gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(KEYINPUT3), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n319), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n326), .A2(new_n250), .A3(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n324), .A2(new_n325), .A3(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT5), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AND2_X1   g131(.A1(new_n312), .A2(new_n319), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(new_n262), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n320), .A2(new_n250), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n325), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n328), .A2(new_n250), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n337), .A2(new_n326), .B1(new_n321), .B2(new_n323), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n336), .B1(new_n338), .B2(new_n325), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n299), .B(new_n332), .C1(new_n339), .C2(new_n331), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT6), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT78), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n299), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n334), .A2(new_n335), .ZN(new_n344));
  INV_X1    g143(.A(new_n325), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n331), .B1(new_n330), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT5), .B1(new_n338), .B2(new_n325), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n343), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n340), .A2(new_n349), .A3(new_n341), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n347), .A2(new_n348), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT78), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT6), .A4(new_n299), .ZN(new_n353));
  AND3_X1   g152(.A1(new_n342), .A2(new_n350), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT72), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  NAND2_X1  g155(.A1(G226gat), .A2(G233gat), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n235), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G211gat), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT69), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT69), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G211gat), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n360), .A2(new_n362), .A3(G218gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT22), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AND2_X1   g164(.A1(G197gat), .A2(G204gat), .ZN(new_n366));
  NOR2_X1   g165(.A1(G197gat), .A2(G204gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  XOR2_X1   g168(.A(G211gat), .B(G218gat), .Z(new_n370));
  AOI22_X1  g169(.A1(new_n365), .A2(new_n369), .B1(KEYINPUT70), .B2(new_n370), .ZN(new_n371));
  OR2_X1    g170(.A1(new_n370), .A2(KEYINPUT70), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  XNOR2_X1  g172(.A(KEYINPUT69), .B(G211gat), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT22), .B1(new_n374), .B2(G218gat), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT71), .ZN(new_n376));
  NOR4_X1   g175(.A1(new_n375), .A2(new_n376), .A3(new_n370), .A4(new_n368), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n368), .B1(new_n363), .B2(new_n364), .ZN(new_n378));
  INV_X1    g177(.A(new_n370), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT71), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n373), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(new_n357), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n223), .B(new_n382), .C1(new_n233), .C2(new_n234), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n358), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n381), .B1(new_n358), .B2(new_n383), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n355), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n365), .A2(new_n379), .A3(new_n369), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n376), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n378), .A2(KEYINPUT71), .A3(new_n379), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n388), .A2(new_n389), .B1(new_n371), .B2(new_n372), .ZN(new_n390));
  NOR3_X1   g189(.A1(new_n261), .A2(KEYINPUT29), .A3(new_n382), .ZN(new_n391));
  INV_X1    g190(.A(new_n383), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n358), .A2(new_n381), .A3(new_n383), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(KEYINPUT72), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n386), .A2(new_n395), .ZN(new_n396));
  XNOR2_X1  g195(.A(KEYINPUT73), .B(G64gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n397), .B(G92gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(G8gat), .B(G36gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n396), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n401), .B1(new_n393), .B2(new_n394), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT30), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT74), .B1(new_n403), .B2(KEYINPUT30), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT74), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT30), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n384), .A2(new_n385), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n406), .B(new_n407), .C1(new_n408), .C2(new_n401), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n402), .A2(new_n404), .A3(new_n405), .A4(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT79), .B1(new_n354), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n342), .A2(new_n350), .A3(new_n353), .ZN(new_n412));
  AND2_X1   g211(.A1(new_n405), .A2(new_n409), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT79), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n396), .A2(new_n401), .B1(KEYINPUT30), .B2(new_n403), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n412), .A2(new_n413), .A3(new_n414), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  XOR2_X1   g216(.A(KEYINPUT31), .B(G50gat), .Z(new_n418));
  XNOR2_X1  g217(.A(G78gat), .B(G106gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT83), .ZN(new_n421));
  INV_X1    g220(.A(G228gat), .ZN(new_n422));
  INV_X1    g221(.A(G233gat), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT80), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n425), .B1(new_n378), .B2(new_n379), .ZN(new_n426));
  OAI211_X1 g225(.A(KEYINPUT80), .B(new_n370), .C1(new_n375), .C2(new_n368), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n388), .A2(new_n389), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT29), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT81), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n327), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n377), .A2(new_n380), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n426), .A2(new_n427), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n356), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n435), .A2(KEYINPUT81), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n320), .B1(new_n432), .B2(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n328), .A2(new_n356), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n381), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n424), .B1(new_n437), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(new_n424), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT82), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n443), .B1(new_n390), .B2(KEYINPUT29), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n381), .A2(KEYINPUT82), .A3(new_n356), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(new_n327), .ZN(new_n446));
  AOI211_X1 g245(.A(new_n442), .B(new_n439), .C1(new_n446), .C2(new_n320), .ZN(new_n447));
  INV_X1    g246(.A(G22gat), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n441), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT3), .B1(new_n435), .B2(KEYINPUT81), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n430), .A2(new_n431), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n333), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n442), .B1(new_n452), .B2(new_n439), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n446), .A2(new_n320), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n454), .A2(new_n424), .A3(new_n440), .ZN(new_n455));
  AOI21_X1  g254(.A(G22gat), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n421), .B1(new_n449), .B2(new_n456), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n448), .B1(new_n441), .B2(new_n447), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n453), .A2(G22gat), .A3(new_n455), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT83), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n453), .A2(new_n460), .A3(new_n455), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n458), .A2(new_n459), .A3(new_n461), .A4(new_n420), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n294), .B1(new_n417), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n342), .A2(new_n353), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT87), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT87), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n342), .A2(new_n468), .A3(new_n353), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NOR3_X1   g269(.A1(new_n384), .A2(new_n385), .A3(new_n355), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT72), .B1(new_n393), .B2(new_n394), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT37), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g272(.A(KEYINPUT86), .B1(new_n408), .B2(KEYINPUT37), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT86), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT37), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n475), .B(new_n476), .C1(new_n384), .C2(new_n385), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n473), .A2(new_n401), .A3(new_n474), .A4(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n403), .B1(new_n478), .B2(KEYINPUT38), .ZN(new_n479));
  AOI21_X1  g278(.A(KEYINPUT38), .B1(new_n408), .B2(KEYINPUT37), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n474), .A2(new_n480), .A3(new_n401), .A4(new_n477), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n470), .A2(new_n479), .A3(new_n350), .A4(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n338), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT39), .ZN(new_n484));
  OR2_X1    g283(.A1(new_n484), .A2(KEYINPUT84), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(KEYINPUT84), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n483), .A2(new_n345), .A3(new_n485), .A4(new_n486), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n344), .A2(new_n345), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT39), .B1(new_n338), .B2(new_n325), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n487), .B(new_n343), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(KEYINPUT40), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n491), .A2(new_n410), .A3(new_n340), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT85), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n491), .A2(new_n410), .A3(KEYINPUT85), .A4(new_n340), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n482), .A2(new_n463), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n286), .B1(new_n282), .B2(new_n283), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(new_n271), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n463), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT35), .B1(new_n500), .B2(new_n417), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n410), .B1(new_n470), .B2(new_n350), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n498), .B1(new_n457), .B2(new_n462), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT35), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI22_X1  g304(.A1(new_n465), .A2(new_n496), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G120gat), .B(G148gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(G176gat), .B(G204gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G230gat), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(new_n423), .ZN(new_n512));
  XNOR2_X1  g311(.A(G57gat), .B(G64gat), .ZN(new_n513));
  INV_X1    g312(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(G71gat), .A2(G78gat), .ZN(new_n515));
  OR2_X1    g314(.A1(G71gat), .A2(G78gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT9), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n515), .B(new_n516), .C1(new_n513), .C2(new_n517), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n520), .A2(KEYINPUT92), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n520), .A2(KEYINPUT92), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524));
  INV_X1    g323(.A(G85gat), .ZN(new_n525));
  INV_X1    g324(.A(G92gat), .ZN(new_n526));
  AOI22_X1  g325(.A1(KEYINPUT8), .A2(new_n524), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT7), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(new_n525), .B2(new_n526), .ZN(new_n529));
  NAND3_X1  g328(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n527), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(G99gat), .B(G106gat), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n531), .B(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n523), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n520), .B(KEYINPUT92), .ZN(new_n535));
  OR2_X1    g334(.A1(new_n531), .A2(new_n532), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n531), .A2(new_n532), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n535), .A2(new_n536), .A3(new_n537), .A4(new_n519), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT10), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n534), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n523), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n541), .A2(KEYINPUT10), .A3(new_n537), .A4(new_n536), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n512), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT99), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  AOI211_X1 g344(.A(KEYINPUT99), .B(new_n512), .C1(new_n540), .C2(new_n542), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n534), .A2(new_n538), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n512), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n510), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n543), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(new_n549), .A3(new_n510), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G15gat), .B(G22gat), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT16), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n556), .B1(new_n557), .B2(G1gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(G1gat), .B2(new_n556), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(G8gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT14), .ZN(new_n562));
  INV_X1    g361(.A(G29gat), .ZN(new_n563));
  INV_X1    g362(.A(G36gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n566));
  AOI22_X1  g365(.A1(new_n565), .A2(new_n566), .B1(G29gat), .B2(G36gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT91), .ZN(new_n568));
  XNOR2_X1  g367(.A(G43gat), .B(G50gat), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n567), .A2(new_n568), .B1(KEYINPUT15), .B2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G43gat), .B(G50gat), .Z(new_n571));
  INV_X1    g370(.A(KEYINPUT15), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(new_n567), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n571), .A2(new_n572), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n567), .B(new_n573), .C1(new_n576), .C2(new_n568), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n575), .A2(KEYINPUT17), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT17), .B1(new_n575), .B2(new_n577), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n561), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n560), .A2(new_n577), .A3(new_n575), .ZN(new_n581));
  NAND2_X1  g380(.A1(G229gat), .A2(G233gat), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT18), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n575), .A2(new_n577), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n561), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(new_n581), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n582), .B(KEYINPUT13), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT18), .A4(new_n582), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n585), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT90), .ZN(new_n593));
  XOR2_X1   g392(.A(G169gat), .B(G197gat), .Z(new_n594));
  XNOR2_X1  g393(.A(G113gat), .B(G141gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XOR2_X1   g395(.A(KEYINPUT88), .B(KEYINPUT11), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(KEYINPUT89), .B(KEYINPUT12), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  AND3_X1   g399(.A1(new_n592), .A2(new_n593), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n600), .B1(new_n592), .B2(new_n593), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NOR3_X1   g403(.A1(new_n506), .A2(new_n555), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT21), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n561), .B(new_n202), .C1(new_n606), .C2(new_n523), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n523), .A2(new_n606), .ZN(new_n608));
  OAI21_X1  g407(.A(G183gat), .B1(new_n608), .B2(new_n560), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(new_n612), .ZN(new_n617));
  AND3_X1   g416(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n541), .A2(KEYINPUT21), .ZN(new_n620));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(new_n359), .ZN(new_n622));
  XNOR2_X1  g421(.A(G127gat), .B(G155gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n620), .B(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n616), .B1(new_n614), .B2(new_n617), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n619), .A2(new_n625), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n625), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(new_n618), .B2(new_n626), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(G232gat), .A2(G233gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT95), .Z(new_n633));
  INV_X1    g432(.A(KEYINPUT41), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g434(.A(G134gat), .B(G162gat), .Z(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT96), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n533), .B1(new_n578), .B2(new_n579), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n633), .A2(new_n634), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  OR2_X1    g441(.A1(new_n586), .A2(new_n533), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n640), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(G190gat), .B(G218gat), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n639), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n640), .A2(new_n645), .A3(new_n642), .A4(new_n643), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n644), .A2(new_n646), .A3(new_n637), .ZN(new_n650));
  INV_X1    g449(.A(new_n639), .ZN(new_n651));
  OR3_X1    g450(.A1(new_n644), .A2(new_n646), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT97), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT97), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n649), .A2(new_n652), .A3(new_n655), .A4(new_n650), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n631), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n658), .A2(KEYINPUT98), .ZN(new_n659));
  INV_X1    g458(.A(KEYINPUT98), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n631), .A2(new_n660), .A3(new_n657), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n605), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n354), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT101), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT100), .B(G1gat), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n666), .B(new_n667), .ZN(G1324gat));
  XOR2_X1   g467(.A(KEYINPUT16), .B(G8gat), .Z(new_n669));
  NAND3_X1  g468(.A1(new_n664), .A2(new_n410), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT42), .ZN(new_n671));
  INV_X1    g470(.A(new_n410), .ZN(new_n672));
  OAI21_X1  g471(.A(G8gat), .B1(new_n663), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n671), .A2(new_n673), .ZN(G1325gat));
  AOI21_X1  g473(.A(G15gat), .B1(new_n664), .B2(new_n499), .ZN(new_n675));
  INV_X1    g474(.A(new_n294), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n663), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n675), .B1(G15gat), .B2(new_n677), .ZN(G1326gat));
  NAND2_X1  g477(.A1(new_n664), .A2(new_n464), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT102), .B(KEYINPUT103), .Z(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g480(.A(KEYINPUT43), .B(G22gat), .Z(new_n682));
  XNOR2_X1  g481(.A(new_n681), .B(new_n682), .ZN(G1327gat));
  INV_X1    g482(.A(KEYINPUT104), .ZN(new_n684));
  OAI21_X1  g483(.A(KEYINPUT44), .B1(new_n506), .B2(new_n657), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n417), .A2(new_n464), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n496), .A2(new_n676), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n501), .A2(new_n505), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  INV_X1    g489(.A(new_n657), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n689), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n631), .A2(new_n604), .A3(new_n555), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n684), .B1(new_n695), .B2(new_n412), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n693), .A2(KEYINPUT104), .A3(new_n354), .A4(new_n694), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(G29gat), .A3(new_n697), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n689), .A2(new_n691), .A3(new_n694), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n699), .A2(new_n563), .A3(new_n354), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n700), .B(KEYINPUT45), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n698), .A2(new_n701), .ZN(G1328gat));
  NAND3_X1  g501(.A1(new_n699), .A2(new_n564), .A3(new_n410), .ZN(new_n703));
  XOR2_X1   g502(.A(new_n703), .B(KEYINPUT46), .Z(new_n704));
  OAI21_X1  g503(.A(G36gat), .B1(new_n695), .B2(new_n672), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1329gat));
  AND3_X1   g505(.A1(new_n699), .A2(new_n273), .A3(new_n499), .ZN(new_n707));
  NAND3_X1  g506(.A1(new_n693), .A2(new_n294), .A3(new_n694), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n707), .B1(G43gat), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g509(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n464), .A2(G50gat), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n699), .A2(new_n464), .ZN(new_n713));
  OAI221_X1 g512(.A(new_n711), .B1(new_n695), .B2(new_n712), .C1(G50gat), .C2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(KEYINPUT105), .A2(KEYINPUT48), .ZN(new_n715));
  XOR2_X1   g514(.A(new_n714), .B(new_n715), .Z(G1331gat));
  NOR2_X1   g515(.A1(new_n506), .A2(new_n554), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n662), .A2(new_n604), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n354), .ZN(new_n721));
  XNOR2_X1  g520(.A(new_n721), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g521(.A1(new_n719), .A2(new_n672), .ZN(new_n723));
  NOR2_X1   g522(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n724));
  AND2_X1   g523(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n723), .B2(new_n724), .ZN(G1333gat));
  OAI21_X1  g526(.A(G71gat), .B1(new_n719), .B2(new_n676), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n720), .A2(new_n499), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n728), .B1(new_n729), .B2(G71gat), .ZN(new_n730));
  XOR2_X1   g529(.A(new_n730), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g530(.A1(new_n720), .A2(new_n464), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G78gat), .ZN(G1335gat));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n631), .A2(new_n603), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n693), .A2(new_n555), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n736), .B2(new_n412), .ZN(new_n737));
  INV_X1    g536(.A(new_n735), .ZN(new_n738));
  AOI211_X1 g537(.A(new_n554), .B(new_n738), .C1(new_n685), .C2(new_n692), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n739), .A2(KEYINPUT106), .A3(new_n354), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n737), .A2(new_n740), .A3(G85gat), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT107), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n506), .B2(new_n657), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n689), .A2(KEYINPUT107), .A3(new_n691), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n743), .A2(new_n744), .A3(new_n735), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT51), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n743), .A2(new_n744), .A3(KEYINPUT51), .A4(new_n735), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n749), .A2(new_n525), .A3(new_n354), .A4(new_n555), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n741), .A2(new_n750), .ZN(G1336gat));
  NOR2_X1   g550(.A1(new_n672), .A2(G92gat), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n749), .A2(new_n555), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n754));
  OAI21_X1  g553(.A(G92gat), .B1(new_n736), .B2(new_n672), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT109), .ZN(new_n757));
  XNOR2_X1  g556(.A(KEYINPUT108), .B(KEYINPUT51), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n745), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n748), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n752), .A2(new_n555), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n755), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n757), .B1(new_n764), .B2(KEYINPUT52), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n526), .B1(new_n739), .B2(new_n410), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n761), .B1(new_n759), .B2(new_n748), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n757), .B(KEYINPUT52), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n756), .B1(new_n765), .B2(new_n769), .ZN(G1337gat));
  OAI21_X1  g569(.A(G99gat), .B1(new_n736), .B2(new_n676), .ZN(new_n771));
  INV_X1    g570(.A(G99gat), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n749), .A2(new_n772), .A3(new_n555), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n773), .B2(new_n498), .ZN(G1338gat));
  NOR3_X1   g573(.A1(new_n463), .A2(G106gat), .A3(new_n554), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n760), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(G106gat), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n777), .B1(new_n739), .B2(new_n464), .ZN(new_n778));
  OAI21_X1  g577(.A(KEYINPUT53), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n749), .A2(new_n775), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT53), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n779), .B1(new_n778), .B2(new_n782), .ZN(G1339gat));
  AND4_X1   g582(.A1(new_n659), .A2(new_n661), .A3(new_n554), .A4(new_n604), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n540), .A2(new_n542), .A3(new_n512), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n543), .B2(KEYINPUT110), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT110), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n540), .A2(new_n542), .A3(new_n787), .A4(new_n512), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(KEYINPUT54), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n545), .B2(new_n546), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n789), .A2(new_n791), .A3(KEYINPUT55), .A4(new_n509), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT111), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n792), .A2(new_n793), .A3(new_n552), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n789), .A2(new_n791), .A3(new_n509), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT55), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n792), .A2(new_n552), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT111), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n585), .A2(new_n590), .A3(new_n591), .A4(new_n600), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n588), .A2(new_n589), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n582), .B1(new_n580), .B2(new_n581), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n598), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n803), .A2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n654), .A2(new_n808), .A3(new_n656), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n799), .A2(new_n800), .A3(new_n802), .A4(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n802), .A2(new_n809), .A3(new_n797), .A4(new_n794), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT112), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n793), .B1(new_n792), .B2(new_n552), .ZN(new_n814));
  NOR3_X1   g613(.A1(new_n798), .A2(new_n604), .A3(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n555), .A2(new_n816), .A3(new_n808), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT113), .B1(new_n554), .B2(new_n807), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n657), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n813), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n631), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n784), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n823), .A2(new_n500), .ZN(new_n824));
  NOR2_X1   g623(.A1(new_n410), .A2(new_n412), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(G113gat), .B1(new_n826), .B2(new_n604), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n603), .A2(new_n238), .ZN(new_n828));
  XOR2_X1   g627(.A(new_n828), .B(KEYINPUT114), .Z(new_n829));
  OAI21_X1  g628(.A(new_n827), .B1(new_n826), .B2(new_n829), .ZN(G1340gat));
  NOR2_X1   g629(.A1(new_n826), .A2(new_n554), .ZN(new_n831));
  XNOR2_X1  g630(.A(KEYINPUT115), .B(G120gat), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n831), .B(new_n832), .ZN(G1341gat));
  NOR2_X1   g632(.A1(new_n826), .A2(new_n822), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(new_n244), .ZN(G1342gat));
  NAND2_X1  g634(.A1(new_n691), .A2(new_n672), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT116), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n824), .A2(new_n242), .A3(new_n354), .A4(new_n838), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n354), .ZN(new_n841));
  OAI21_X1  g640(.A(G134gat), .B1(new_n841), .B2(new_n836), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n840), .A2(new_n842), .A3(new_n843), .ZN(G1343gat));
  NAND2_X1  g643(.A1(new_n676), .A2(new_n825), .ZN(new_n845));
  XNOR2_X1  g644(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n795), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n792), .A2(new_n552), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n795), .A2(KEYINPUT118), .A3(new_n846), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n849), .A2(new_n850), .A3(new_n603), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n555), .A2(new_n808), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT119), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(KEYINPUT119), .A3(new_n853), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n856), .A2(new_n657), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n631), .B1(new_n858), .B2(new_n813), .ZN(new_n859));
  OAI211_X1 g658(.A(KEYINPUT57), .B(new_n464), .C1(new_n859), .C2(new_n784), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT57), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n861), .B1(new_n823), .B2(new_n463), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n845), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n863), .A2(G141gat), .A3(new_n603), .ZN(new_n864));
  INV_X1    g663(.A(new_n823), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n294), .A2(KEYINPUT120), .A3(new_n463), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n412), .ZN(new_n867));
  OAI21_X1  g666(.A(KEYINPUT120), .B1(new_n294), .B2(new_n463), .ZN(new_n868));
  NAND4_X1  g667(.A1(new_n865), .A2(new_n672), .A3(new_n867), .A4(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n302), .B1(new_n869), .B2(new_n604), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n864), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n871), .B(new_n872), .ZN(G1344gat));
  AOI21_X1  g672(.A(new_n631), .B1(new_n858), .B2(new_n811), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n861), .B(new_n464), .C1(new_n874), .C2(new_n784), .ZN(new_n875));
  OAI21_X1  g674(.A(KEYINPUT57), .B1(new_n823), .B2(new_n463), .ZN(new_n876));
  INV_X1    g675(.A(new_n845), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n555), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(G148gat), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT59), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n860), .A2(new_n862), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n881), .A2(new_n555), .A3(new_n877), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n304), .A2(KEYINPUT59), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n882), .A2(KEYINPUT121), .A3(new_n883), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT121), .B1(new_n882), .B2(new_n883), .ZN(new_n885));
  OAI21_X1  g684(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(new_n869), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n304), .A3(new_n555), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n886), .A2(new_n888), .ZN(G1345gat));
  AOI21_X1  g688(.A(G155gat), .B1(new_n887), .B2(new_n631), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n822), .A2(new_n309), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n890), .B1(new_n863), .B2(new_n891), .ZN(G1346gat));
  NOR2_X1   g691(.A1(new_n837), .A2(G162gat), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n865), .A2(new_n867), .A3(new_n868), .A4(new_n893), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n863), .A2(new_n691), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n894), .B1(new_n895), .B2(new_n310), .ZN(G1347gat));
  NOR2_X1   g695(.A1(new_n672), .A2(new_n354), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n631), .B1(new_n813), .B2(new_n820), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n503), .B(new_n897), .C1(new_n898), .C2(new_n784), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT122), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n899), .B(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(G169gat), .B1(new_n901), .B2(new_n604), .ZN(new_n902));
  INV_X1    g701(.A(new_n899), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n214), .A3(new_n603), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1348gat));
  OAI21_X1  g704(.A(G176gat), .B1(new_n901), .B2(new_n554), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n899), .A2(G176gat), .A3(new_n554), .ZN(new_n908));
  INV_X1    g707(.A(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n907), .B1(new_n906), .B2(new_n909), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(G1349gat));
  INV_X1    g712(.A(KEYINPUT124), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n631), .A2(new_n211), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n899), .B2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n822), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n202), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT60), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n921), .B(new_n917), .C1(new_n918), .C2(new_n202), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1350gat));
  NAND3_X1  g722(.A1(new_n903), .A2(new_n207), .A3(new_n691), .ZN(new_n924));
  XNOR2_X1  g723(.A(new_n899), .B(KEYINPUT122), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n207), .B1(new_n925), .B2(new_n691), .ZN(new_n926));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n927));
  AND2_X1   g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n924), .B1(new_n928), .B2(new_n929), .ZN(G1351gat));
  XOR2_X1   g729(.A(KEYINPUT126), .B(G197gat), .Z(new_n931));
  AND2_X1   g730(.A1(new_n875), .A2(new_n876), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n676), .A2(new_n897), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n931), .B1(new_n935), .B2(new_n604), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n865), .A2(new_n464), .A3(new_n934), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT125), .ZN(new_n938));
  XNOR2_X1  g737(.A(new_n937), .B(new_n938), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n939), .A2(new_n931), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n936), .B1(new_n940), .B2(new_n604), .ZN(G1352gat));
  NOR3_X1   g740(.A1(new_n937), .A2(G204gat), .A3(new_n554), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  NOR4_X1   g744(.A1(new_n937), .A2(KEYINPUT127), .A3(G204gat), .A4(new_n554), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n945), .A2(KEYINPUT62), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n932), .A2(new_n555), .A3(new_n934), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G204gat), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT62), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n951), .B1(new_n944), .B2(new_n946), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n948), .A2(new_n950), .A3(new_n952), .ZN(G1353gat));
  NAND3_X1  g752(.A1(new_n932), .A2(new_n631), .A3(new_n934), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n954), .B2(G211gat), .ZN(new_n956));
  OR2_X1    g755(.A1(new_n822), .A2(new_n374), .ZN(new_n957));
  OAI22_X1  g756(.A1(new_n955), .A2(new_n956), .B1(new_n939), .B2(new_n957), .ZN(G1354gat));
  OAI21_X1  g757(.A(G218gat), .B1(new_n935), .B2(new_n657), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n939), .A2(G218gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n959), .B1(new_n960), .B2(new_n657), .ZN(G1355gat));
endmodule


