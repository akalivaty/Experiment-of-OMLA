//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n539,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n569, new_n570, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n586, new_n587, new_n589, new_n590,
    new_n591, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n630, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  XOR2_X1   g026(.A(KEYINPUT64), .B(KEYINPUT65), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n451), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n451), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n461), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(KEYINPUT66), .A3(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n467));
  NAND4_X1  g042(.A1(new_n463), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G137), .ZN(new_n469));
  INV_X1    g044(.A(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n466), .A2(G2104), .ZN(new_n471));
  OAI22_X1  g046(.A1(new_n468), .A2(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT67), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n474));
  OAI221_X1 g049(.A(new_n474), .B1(new_n470), .B2(new_n471), .C1(new_n468), .C2(new_n469), .ZN(new_n475));
  AND2_X1   g050(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(G113), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n464), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n467), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G125), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  OAI21_X1  g059(.A(KEYINPUT68), .B1(G100), .B2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  NOR3_X1   g061(.A1(KEYINPUT68), .A2(G100), .A3(G2105), .ZN(new_n487));
  OAI221_X1 g062(.A(G2104), .B1(G112), .B2(new_n466), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n463), .A2(new_n467), .A3(new_n465), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n489), .A2(new_n466), .ZN(new_n490));
  INV_X1    g065(.A(G124), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(new_n468), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n492), .B1(G136), .B2(new_n493), .ZN(new_n494));
  XOR2_X1   g069(.A(new_n494), .B(KEYINPUT69), .Z(G162));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n463), .A2(new_n465), .A3(new_n497), .A4(new_n467), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(KEYINPUT4), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n467), .A2(new_n478), .ZN(new_n500));
  NOR3_X1   g075(.A1(new_n496), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  AND2_X1   g078(.A1(G126), .A2(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n463), .A2(new_n465), .A3(new_n467), .A4(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n466), .A2(G114), .ZN(new_n507));
  OAI21_X1  g082(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OR2_X1    g084(.A1(G102), .A2(G2105), .ZN(new_n510));
  INV_X1    g085(.A(G114), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G2105), .ZN(new_n512));
  NAND4_X1  g087(.A1(new_n510), .A2(new_n512), .A3(KEYINPUT70), .A4(G2104), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n503), .A2(new_n505), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  OR2_X1    g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI22_X1  g094(.A1(new_n519), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n520));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT6), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n524), .B2(new_n521), .ZN(new_n525));
  NAND3_X1  g100(.A1(KEYINPUT71), .A2(KEYINPUT6), .A3(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(new_n519), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(G88), .ZN(new_n530));
  INV_X1    g105(.A(G543), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n531), .B1(new_n525), .B2(new_n526), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(G50), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT72), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n530), .A2(new_n536), .A3(new_n533), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n522), .B1(new_n535), .B2(new_n537), .ZN(G166));
  NAND3_X1  g113(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT73), .ZN(new_n540));
  NAND3_X1  g115(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n541), .A2(KEYINPUT7), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n532), .A2(G51), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n529), .A2(G89), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n540), .A2(new_n544), .A3(new_n545), .ZN(G286));
  INV_X1    g121(.A(G286), .ZN(G168));
  NAND2_X1  g122(.A1(new_n529), .A2(G90), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n532), .A2(G52), .ZN(new_n549));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  XOR2_X1   g125(.A(KEYINPUT5), .B(G543), .Z(new_n551));
  INV_X1    g126(.A(G64), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  AND4_X1   g129(.A1(KEYINPUT74), .A2(new_n548), .A3(new_n549), .A4(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n529), .A2(G90), .B1(new_n553), .B2(G651), .ZN(new_n556));
  AOI21_X1  g131(.A(KEYINPUT74), .B1(new_n556), .B2(new_n549), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n555), .A2(new_n557), .ZN(G301));
  INV_X1    g133(.A(G301), .ZN(G171));
  NAND2_X1  g134(.A1(G68), .A2(G543), .ZN(new_n560));
  INV_X1    g135(.A(G56), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n551), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n529), .A2(G81), .B1(new_n562), .B2(G651), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n532), .A2(G43), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  AND2_X1   g146(.A1(KEYINPUT75), .A2(G53), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n532), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(KEYINPUT9), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT9), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n532), .A2(new_n575), .A3(new_n572), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n574), .A2(new_n576), .B1(G91), .B2(new_n529), .ZN(new_n577));
  INV_X1    g152(.A(G65), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n551), .A2(KEYINPUT76), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n519), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n578), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g157(.A1(G78), .A2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n577), .A2(new_n584), .ZN(G299));
  NAND2_X1  g160(.A1(new_n535), .A2(new_n537), .ZN(new_n586));
  INV_X1    g161(.A(new_n522), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G303));
  NAND2_X1  g163(.A1(new_n529), .A2(G87), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n532), .A2(G49), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n519), .B2(G74), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(G288));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(KEYINPUT77), .B1(new_n551), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n519), .A2(new_n595), .A3(G61), .ZN(new_n596));
  NAND2_X1  g171(.A1(G73), .A2(G543), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n594), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(G86), .B2(new_n529), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n532), .A2(G48), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT78), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n599), .A2(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n532), .A2(G47), .ZN(new_n603));
  INV_X1    g178(.A(G85), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n605));
  OAI221_X1 g180(.A(new_n603), .B1(new_n528), .B2(new_n604), .C1(new_n521), .C2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT79), .ZN(G290));
  INV_X1    g182(.A(G868), .ZN(new_n608));
  NOR2_X1   g183(.A1(G301), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n529), .A2(KEYINPUT10), .A3(G92), .ZN(new_n610));
  INV_X1    g185(.A(KEYINPUT10), .ZN(new_n611));
  INV_X1    g186(.A(G92), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n528), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT80), .B(G66), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n615), .B1(new_n579), .B2(new_n581), .ZN(new_n616));
  AND2_X1   g191(.A1(G79), .A2(G543), .ZN(new_n617));
  OAI21_X1  g192(.A(G651), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n532), .A2(G54), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n614), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AND2_X1   g195(.A1(new_n620), .A2(KEYINPUT81), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n620), .A2(KEYINPUT81), .ZN(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n609), .B1(new_n623), .B2(new_n608), .ZN(G284));
  AOI21_X1  g199(.A(new_n609), .B1(new_n623), .B2(new_n608), .ZN(G321));
  NAND2_X1  g200(.A1(G286), .A2(G868), .ZN(new_n626));
  INV_X1    g201(.A(G299), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G868), .ZN(G280));
  XNOR2_X1  g203(.A(G280), .B(KEYINPUT82), .ZN(G297));
  XOR2_X1   g204(.A(KEYINPUT83), .B(G559), .Z(new_n630));
  OAI21_X1  g205(.A(new_n623), .B1(G860), .B2(new_n630), .ZN(G148));
  NAND2_X1  g206(.A1(new_n565), .A2(new_n608), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n623), .A2(new_n630), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n632), .B1(new_n634), .B2(new_n608), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g211(.A(new_n471), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n500), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  INV_X1    g216(.A(G123), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n643));
  NOR3_X1   g218(.A1(new_n643), .A2(new_n466), .A3(G111), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n643), .B1(new_n466), .B2(G111), .ZN(new_n645));
  OR2_X1    g220(.A1(G99), .A2(G2105), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(G2104), .A3(new_n646), .ZN(new_n647));
  OAI22_X1  g222(.A1(new_n490), .A2(new_n642), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(G135), .B2(new_n493), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n650), .A2(G2096), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(G2096), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n641), .A2(new_n651), .A3(new_n652), .ZN(G156));
  XNOR2_X1  g228(.A(G2427), .B(G2438), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2430), .ZN(new_n655));
  XNOR2_X1  g230(.A(KEYINPUT15), .B(G2435), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n656), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(KEYINPUT14), .A3(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G1341), .B(G1348), .Z(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n659), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(KEYINPUT85), .B(KEYINPUT16), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n664), .B(new_n665), .Z(new_n666));
  OR2_X1    g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n663), .A2(new_n666), .ZN(new_n668));
  AND3_X1   g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(G401));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  XNOR2_X1  g246(.A(G2067), .B(G2678), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n670), .B1(new_n673), .B2(KEYINPUT18), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT86), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G2100), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT18), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n673), .A2(KEYINPUT17), .ZN(new_n678));
  NOR2_X1   g253(.A1(new_n671), .A2(new_n672), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(G2096), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n676), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT20), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n685), .A2(new_n686), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n684), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n684), .B2(new_n690), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G229));
  NAND3_X1  g274(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT90), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n701), .A2(KEYINPUT25), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(KEYINPUT25), .ZN(new_n703));
  NAND2_X1  g278(.A1(G115), .A2(G2104), .ZN(new_n704));
  INV_X1    g279(.A(G127), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n479), .B2(new_n705), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n702), .A2(new_n703), .B1(G2105), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n493), .A2(G139), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT91), .Z(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n711), .B2(G33), .ZN(new_n713));
  INV_X1    g288(.A(G2072), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT24), .B(G34), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(new_n711), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT92), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n483), .B2(new_n711), .ZN(new_n719));
  INV_X1    g294(.A(G2084), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G20), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT23), .Z(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(G299), .B2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G1956), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NOR4_X1   g303(.A1(new_n715), .A2(new_n721), .A3(new_n722), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n723), .A2(G5), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G171), .B2(new_n723), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n731), .A2(G1961), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT95), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n723), .A2(G4), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n623), .B2(new_n723), .ZN(new_n735));
  AND2_X1   g310(.A1(new_n735), .A2(G1348), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n735), .A2(G1348), .ZN(new_n737));
  NOR3_X1   g312(.A1(new_n733), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n711), .A2(G32), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT26), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n740), .A2(new_n741), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n742), .A2(new_n743), .B1(G105), .B2(new_n637), .ZN(new_n744));
  INV_X1    g319(.A(G129), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n490), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G141), .B2(new_n493), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(new_n711), .ZN(new_n748));
  XNOR2_X1  g323(.A(KEYINPUT27), .B(G1996), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NOR2_X1   g325(.A1(G164), .A2(new_n711), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G27), .B2(new_n711), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n752), .A2(new_n753), .ZN(new_n755));
  NAND3_X1  g330(.A1(new_n750), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n711), .A2(G26), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT28), .ZN(new_n758));
  OR2_X1    g333(.A1(G104), .A2(G2105), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n759), .B(G2104), .C1(G116), .C2(new_n466), .ZN(new_n760));
  INV_X1    g335(.A(G128), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n490), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G140), .B2(new_n493), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n758), .B1(new_n763), .B2(new_n711), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT89), .ZN(new_n765));
  INV_X1    g340(.A(G2067), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n756), .B(new_n767), .C1(new_n713), .C2(new_n714), .ZN(new_n768));
  NOR2_X1   g343(.A1(G168), .A2(new_n723), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n723), .B2(G21), .ZN(new_n770));
  XNOR2_X1  g345(.A(KEYINPUT93), .B(G1966), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT94), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n711), .A2(G35), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G162), .B2(new_n711), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT29), .B(G2090), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n775), .B(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n731), .A2(G1961), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n723), .A2(G19), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n566), .B2(new_n723), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(G1341), .Z(new_n781));
  INV_X1    g356(.A(G11), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n782), .A2(KEYINPUT31), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(KEYINPUT31), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT30), .ZN(new_n785));
  AND2_X1   g360(.A1(new_n785), .A2(G28), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n711), .B1(new_n785), .B2(G28), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n783), .B(new_n784), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n649), .B2(G29), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n781), .B(new_n789), .C1(new_n770), .C2(new_n771), .ZN(new_n790));
  NOR4_X1   g365(.A1(new_n773), .A2(new_n777), .A3(new_n778), .A4(new_n790), .ZN(new_n791));
  NAND4_X1  g366(.A1(new_n729), .A2(new_n738), .A3(new_n768), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n723), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n723), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1971), .ZN(new_n795));
  INV_X1    g370(.A(KEYINPUT88), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n795), .A2(new_n796), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n723), .A2(G23), .ZN(new_n799));
  INV_X1    g374(.A(G288), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n799), .B1(new_n800), .B2(new_n723), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT87), .ZN(new_n802));
  XOR2_X1   g377(.A(KEYINPUT33), .B(G1976), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n802), .B(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(G6), .A2(G16), .ZN(new_n805));
  INV_X1    g380(.A(G305), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n805), .B1(new_n806), .B2(G16), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT32), .B(G1981), .Z(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  AND4_X1   g384(.A1(new_n797), .A2(new_n798), .A3(new_n804), .A4(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT34), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n711), .A2(G25), .ZN(new_n814));
  INV_X1    g389(.A(G119), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n466), .A2(G107), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n817));
  OAI22_X1  g392(.A1(new_n490), .A2(new_n815), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n493), .A2(G131), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n814), .B1(new_n820), .B2(new_n711), .ZN(new_n821));
  XNOR2_X1  g396(.A(KEYINPUT35), .B(G1991), .ZN(new_n822));
  XOR2_X1   g397(.A(new_n821), .B(new_n822), .Z(new_n823));
  INV_X1    g398(.A(G290), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(new_n723), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n723), .B2(G24), .ZN(new_n826));
  INV_X1    g401(.A(G1986), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n827), .B2(new_n826), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n812), .A2(new_n813), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n831));
  AND2_X1   g406(.A1(new_n813), .A2(new_n829), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT36), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n832), .A2(new_n833), .A3(new_n812), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n792), .B1(new_n831), .B2(new_n834), .ZN(G311));
  INV_X1    g410(.A(new_n792), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n833), .B1(new_n832), .B2(new_n812), .ZN(new_n837));
  AND4_X1   g412(.A1(new_n833), .A2(new_n812), .A3(new_n813), .A4(new_n829), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n836), .B1(new_n837), .B2(new_n838), .ZN(G150));
  NAND2_X1  g414(.A1(G80), .A2(G543), .ZN(new_n840));
  INV_X1    g415(.A(G67), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n551), .B2(new_n841), .ZN(new_n842));
  AOI22_X1  g417(.A1(new_n529), .A2(G93), .B1(new_n842), .B2(G651), .ZN(new_n843));
  XNOR2_X1  g418(.A(KEYINPUT97), .B(G55), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n532), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(G860), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT99), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT37), .ZN(new_n849));
  INV_X1    g424(.A(G860), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n623), .A2(G559), .ZN(new_n851));
  XOR2_X1   g426(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n851), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n565), .A2(new_n846), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n563), .A2(new_n843), .A3(new_n564), .A4(new_n845), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n851), .B(new_n852), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n860), .A2(new_n857), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n850), .B1(new_n862), .B2(KEYINPUT39), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT98), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(KEYINPUT39), .ZN(new_n866));
  AND3_X1   g441(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n865), .B1(new_n864), .B2(new_n866), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n849), .B1(new_n867), .B2(new_n868), .ZN(G145));
  XNOR2_X1  g444(.A(new_n483), .B(new_n649), .ZN(new_n870));
  XNOR2_X1  g445(.A(G162), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT100), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n514), .A2(new_n872), .A3(new_n505), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n872), .B1(new_n514), .B2(new_n505), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n503), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n763), .B(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(new_n747), .ZN(new_n877));
  INV_X1    g452(.A(new_n709), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n710), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n880), .B2(new_n877), .ZN(new_n881));
  OAI21_X1  g456(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n882));
  INV_X1    g457(.A(G118), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n882), .B1(new_n883), .B2(G2105), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n493), .A2(G142), .ZN(new_n885));
  XOR2_X1   g460(.A(new_n885), .B(KEYINPUT101), .Z(new_n886));
  INV_X1    g461(.A(new_n490), .ZN(new_n887));
  AOI211_X1 g462(.A(new_n884), .B(new_n886), .C1(G130), .C2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n820), .B(new_n639), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n881), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n881), .A2(new_n890), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n871), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n893), .ZN(new_n895));
  INV_X1    g470(.A(new_n871), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n896), .A3(new_n891), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n894), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g475(.A(new_n633), .B(new_n858), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT41), .ZN(new_n902));
  NAND2_X1  g477(.A1(G299), .A2(KEYINPUT102), .ZN(new_n903));
  INV_X1    g478(.A(new_n620), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT102), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n577), .A2(new_n905), .A3(new_n584), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n620), .A2(G299), .A3(KEYINPUT102), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n902), .B1(new_n907), .B2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n903), .A2(new_n904), .A3(new_n906), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n911), .A2(KEYINPUT41), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n901), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n907), .A2(new_n909), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n914), .B1(new_n901), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT42), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n914), .B(new_n918), .C1(new_n901), .C2(new_n915), .ZN(new_n919));
  NAND2_X1  g494(.A1(G290), .A2(G166), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n824), .A2(G303), .ZN(new_n921));
  XNOR2_X1  g496(.A(G288), .B(KEYINPUT103), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(G305), .ZN(new_n923));
  OR2_X1    g498(.A1(new_n922), .A2(G305), .ZN(new_n924));
  AND4_X1   g499(.A1(new_n920), .A2(new_n921), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  AOI22_X1  g500(.A1(new_n923), .A2(new_n924), .B1(new_n921), .B2(new_n920), .ZN(new_n926));
  NOR2_X1   g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n927), .A2(KEYINPUT104), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n917), .A2(new_n919), .A3(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n928), .B1(new_n917), .B2(new_n919), .ZN(new_n930));
  OAI21_X1  g505(.A(G868), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n846), .A2(new_n608), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n931), .A2(new_n932), .ZN(G295));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n932), .ZN(G331));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(new_n555), .B2(new_n557), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n548), .A2(new_n549), .A3(new_n554), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT74), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n556), .A2(KEYINPUT74), .A3(new_n549), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT105), .ZN(new_n942));
  AND3_X1   g517(.A1(new_n937), .A2(new_n857), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n857), .B1(new_n937), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g519(.A(G286), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n937), .A2(new_n942), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n858), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n937), .A2(new_n857), .A3(new_n942), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(G168), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n945), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n912), .ZN(new_n951));
  AOI21_X1  g526(.A(KEYINPUT41), .B1(new_n911), .B2(new_n908), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n945), .A2(new_n949), .A3(new_n915), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n925), .A2(new_n926), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT106), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n945), .A2(new_n949), .A3(KEYINPUT106), .A4(new_n915), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n960), .A2(new_n954), .A3(new_n927), .A4(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT43), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n958), .A2(new_n962), .A3(new_n963), .A4(new_n898), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT107), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n962), .A2(new_n898), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n955), .A2(new_n959), .B1(new_n950), .B2(new_n953), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n927), .B1(new_n968), .B2(new_n961), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT43), .B1(new_n967), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n964), .A2(new_n965), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n935), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n963), .B1(new_n967), .B2(new_n969), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n958), .A2(new_n962), .A3(new_n898), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(new_n975), .B2(new_n963), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT44), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n973), .A2(new_n977), .ZN(G397));
  INV_X1    g553(.A(KEYINPUT51), .ZN(new_n979));
  INV_X1    g554(.A(G8), .ZN(new_n980));
  INV_X1    g555(.A(G40), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(new_n481), .B2(G2105), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n473), .A2(new_n475), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT50), .B1(new_n875), .B2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n515), .A2(KEYINPUT50), .A3(new_n984), .ZN(new_n986));
  INV_X1    g561(.A(new_n986), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n720), .B(new_n983), .C1(new_n985), .C2(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT45), .B1(new_n875), .B2(new_n984), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT45), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n990), .A2(G1384), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n515), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n983), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n771), .B1(new_n989), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n980), .B1(new_n988), .B2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n979), .B1(new_n995), .B2(G286), .ZN(new_n996));
  NAND2_X1  g571(.A1(G286), .A2(G8), .ZN(new_n997));
  XOR2_X1   g572(.A(new_n997), .B(KEYINPUT119), .Z(new_n998));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n998), .B1(new_n995), .B2(new_n999), .ZN(new_n1000));
  AOI211_X1 g575(.A(KEYINPUT118), .B(new_n980), .C1(new_n988), .C2(new_n994), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n996), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT120), .ZN(new_n1003));
  INV_X1    g578(.A(new_n995), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(new_n979), .A3(new_n997), .ZN(new_n1005));
  AND3_X1   g580(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1003), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1007));
  OAI21_X1  g582(.A(KEYINPUT62), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1002), .A2(new_n1005), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT120), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT62), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(G1981), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n1014), .B1(new_n599), .B2(new_n601), .ZN(new_n1015));
  INV_X1    g590(.A(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n599), .A2(new_n601), .A3(new_n1014), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT114), .ZN(new_n1018));
  OAI211_X1 g593(.A(new_n1016), .B(new_n1017), .C1(new_n1018), .C2(KEYINPUT49), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n983), .A2(new_n984), .A3(new_n875), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(new_n980), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1018), .A2(KEYINPUT49), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1017), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1023), .B1(new_n1024), .B2(new_n1015), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1019), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n800), .A2(G1976), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1020), .A2(new_n1027), .A3(G8), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n800), .A2(G1976), .ZN(new_n1029));
  OR3_X1    g604(.A1(new_n1028), .A2(KEYINPUT52), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(KEYINPUT52), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1026), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1033), .B1(new_n875), .B2(new_n984), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n514), .A2(new_n505), .ZN(new_n1036));
  AOI22_X1  g611(.A1(new_n498), .A2(KEYINPUT4), .B1(new_n500), .B2(new_n501), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1033), .B(new_n984), .C1(new_n1036), .C2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n983), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G2090), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1035), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n984), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n990), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1036), .A2(KEYINPUT100), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n514), .A2(new_n872), .A3(new_n505), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1037), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n991), .ZN(new_n1048));
  OAI211_X1 g623(.A(new_n983), .B(new_n1044), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT110), .B(G1971), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n980), .B1(new_n1042), .B2(new_n1051), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT113), .B(KEYINPUT55), .ZN(new_n1053));
  NAND3_X1  g628(.A1(G303), .A2(G8), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1053), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(G166), .B2(new_n980), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1052), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1032), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT112), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT111), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1049), .A2(new_n1061), .A3(new_n1050), .ZN(new_n1062));
  OAI211_X1 g637(.A(new_n1041), .B(new_n983), .C1(new_n985), .C2(new_n987), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1061), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1060), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1065), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1067), .A2(KEYINPUT112), .A3(new_n1062), .A4(new_n1063), .ZN(new_n1068));
  NAND4_X1  g643(.A1(new_n1066), .A2(new_n1068), .A3(G8), .A4(new_n1057), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1059), .A2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n983), .B1(new_n985), .B2(new_n987), .ZN(new_n1071));
  INV_X1    g646(.A(G1961), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n989), .A2(new_n993), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(KEYINPUT53), .A3(new_n753), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1076), .B1(new_n1049), .B2(G2078), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1073), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1078), .A2(new_n1079), .A3(G171), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(G171), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(KEYINPUT121), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1070), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1008), .A2(new_n1013), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n1086));
  AND3_X1   g661(.A1(new_n577), .A2(new_n1086), .A3(new_n584), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1086), .B1(new_n577), .B2(new_n584), .ZN(new_n1088));
  NOR2_X1   g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n727), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n875), .A2(new_n991), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT56), .B(G2072), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1091), .A2(new_n983), .A3(new_n1044), .A4(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1089), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G1348), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1071), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n983), .A2(new_n984), .A3(new_n875), .A4(new_n766), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n1097), .B(KEYINPUT116), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n623), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1090), .A2(new_n1089), .A3(new_n1093), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1094), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT117), .B(KEYINPUT60), .Z(new_n1103));
  INV_X1    g678(.A(KEYINPUT60), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n1097), .B(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1071), .A2(new_n1095), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI211_X1 g683(.A(new_n1099), .B(new_n1103), .C1(new_n1108), .C2(new_n623), .ZN(new_n1109));
  XNOR2_X1  g684(.A(KEYINPUT58), .B(G1341), .ZN(new_n1110));
  OAI22_X1  g685(.A1(new_n1021), .A2(new_n1110), .B1(new_n1049), .B2(G1996), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n566), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT59), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1101), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT61), .B1(new_n1114), .B2(new_n1094), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1089), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT61), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1118), .A2(new_n1119), .A3(new_n1101), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1115), .A2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1109), .A2(new_n1113), .A3(new_n1121), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT60), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1123));
  INV_X1    g698(.A(new_n623), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1103), .B1(new_n1125), .B2(new_n1099), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1102), .B1(new_n1122), .B2(new_n1126), .ZN(new_n1127));
  AND2_X1   g702(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n983), .B(KEYINPUT122), .ZN(new_n1129));
  INV_X1    g704(.A(new_n989), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1076), .B1(KEYINPUT123), .B2(new_n753), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(KEYINPUT123), .B2(new_n753), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1132), .B1(new_n875), .B2(new_n991), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1129), .A2(new_n1130), .A3(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1128), .A2(KEYINPUT124), .A3(G301), .A4(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT124), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1073), .A3(new_n1077), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1136), .B1(new_n1137), .B2(G171), .ZN(new_n1138));
  NAND4_X1  g713(.A1(new_n1082), .A2(new_n1135), .A3(new_n1138), .A4(new_n1080), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT54), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1070), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1128), .A2(G301), .A3(new_n1075), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1137), .A2(G171), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(new_n1143), .A3(KEYINPUT54), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1144), .A2(KEYINPUT125), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1142), .A2(new_n1143), .A3(new_n1146), .A4(KEYINPUT54), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1145), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1085), .A2(new_n1127), .A3(new_n1141), .A4(new_n1148), .ZN(new_n1149));
  NOR2_X1   g724(.A1(G288), .A2(G1976), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1024), .B1(new_n1026), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(KEYINPUT115), .ZN(new_n1152));
  AND2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1022), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1154));
  OAI22_X1  g729(.A1(new_n1153), .A2(new_n1154), .B1(new_n1069), .B2(new_n1032), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT63), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n995), .A2(G168), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1156), .B1(new_n1070), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1066), .A2(new_n1068), .A3(G8), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1159), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1032), .A2(new_n1157), .A3(new_n1156), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1160), .A2(new_n1069), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1155), .B1(new_n1158), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1084), .A2(new_n1149), .A3(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n989), .A2(new_n983), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n763), .B(G2067), .ZN(new_n1166));
  INV_X1    g741(.A(G1996), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n747), .A2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1165), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1165), .A2(new_n1167), .A3(new_n747), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT109), .ZN(new_n1171));
  OR2_X1    g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1169), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n820), .B(new_n822), .Z(new_n1175));
  INV_X1    g750(.A(new_n1165), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AND2_X1   g752(.A1(new_n1174), .A2(new_n1177), .ZN(new_n1178));
  NOR3_X1   g753(.A1(new_n824), .A2(new_n1165), .A3(new_n827), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1165), .A2(G290), .A3(G1986), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  XOR2_X1   g756(.A(new_n1181), .B(KEYINPUT108), .Z(new_n1182));
  AND2_X1   g757(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1164), .A2(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT46), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n1165), .B2(G1996), .ZN(new_n1186));
  XOR2_X1   g761(.A(new_n1186), .B(KEYINPUT126), .Z(new_n1187));
  OAI211_X1 g762(.A(new_n1166), .B(new_n747), .C1(new_n1185), .C2(G1996), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1188), .A2(new_n1176), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1187), .A2(new_n1189), .ZN(new_n1190));
  XNOR2_X1  g765(.A(new_n1190), .B(KEYINPUT47), .ZN(new_n1191));
  OR2_X1    g766(.A1(new_n1191), .A2(KEYINPUT127), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1191), .A2(KEYINPUT127), .ZN(new_n1193));
  NOR3_X1   g768(.A1(new_n818), .A2(new_n822), .A3(new_n819), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1174), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n763), .A2(new_n766), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1165), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1180), .B(KEYINPUT48), .Z(new_n1198));
  AOI21_X1  g773(.A(new_n1197), .B1(new_n1178), .B2(new_n1198), .ZN(new_n1199));
  AND3_X1   g774(.A1(new_n1192), .A2(new_n1193), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1184), .A2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g776(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1203));
  OAI211_X1 g777(.A(new_n899), .B(new_n1203), .C1(new_n971), .C2(new_n972), .ZN(G225));
  INV_X1    g778(.A(G225), .ZN(G308));
endmodule


