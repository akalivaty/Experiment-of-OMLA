//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:57 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n570, new_n572, new_n573,
    new_n574, new_n576, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n624, new_n626,
    new_n627, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT66), .B(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT67), .B(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT68), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT69), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  AND3_X1   g044(.A1(new_n463), .A2(new_n465), .A3(new_n469), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n468), .A2(G2105), .B1(G137), .B2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT70), .B1(new_n462), .B2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT70), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(new_n469), .A3(G2104), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G101), .ZN(new_n476));
  OAI21_X1  g051(.A(KEYINPUT71), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT71), .ZN(new_n478));
  NAND4_X1  g053(.A1(new_n472), .A2(new_n474), .A3(new_n478), .A4(G101), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n471), .A2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n466), .A2(new_n469), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n470), .A2(G136), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n483), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NAND2_X1  g063(.A1(new_n469), .A2(G2104), .ZN(new_n489));
  INV_X1    g064(.A(G102), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n463), .A2(new_n465), .A3(G126), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n491), .B1(new_n494), .B2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G138), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n497), .A2(new_n463), .A3(new_n465), .A4(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT72), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT3), .B(G2104), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT73), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n504), .A2(new_n501), .A3(new_n497), .A4(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n495), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  AND2_X1   g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT75), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n515), .A2(new_n516), .A3(G62), .ZN(new_n517));
  NAND2_X1  g092(.A1(G75), .A2(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n512), .A2(new_n514), .ZN(new_n519));
  INV_X1    g094(.A(G62), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT75), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n517), .A2(new_n518), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT74), .A2(G651), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(KEYINPUT74), .A2(KEYINPUT6), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n527), .ZN(new_n531));
  AOI21_X1  g106(.A(KEYINPUT6), .B1(KEYINPUT74), .B2(G651), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n519), .ZN(new_n534));
  AOI22_X1  g109(.A1(G50), .A2(new_n530), .B1(new_n534), .B2(G88), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n523), .A2(new_n535), .ZN(G303));
  INV_X1    g111(.A(G303), .ZN(G166));
  NAND3_X1  g112(.A1(new_n515), .A2(G63), .A3(G651), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT76), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n538), .B(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT77), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n529), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g117(.A1(new_n528), .A2(KEYINPUT77), .A3(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G51), .ZN(new_n545));
  NAND3_X1  g120(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n546));
  XOR2_X1   g121(.A(new_n546), .B(KEYINPUT7), .Z(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n534), .B2(G89), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n540), .A2(new_n545), .A3(new_n548), .ZN(G286));
  INV_X1    g124(.A(G286), .ZN(G168));
  NAND2_X1  g125(.A1(G77), .A2(G543), .ZN(new_n551));
  INV_X1    g126(.A(G64), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n519), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  INV_X1    g129(.A(G90), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n515), .A2(new_n528), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n557), .B1(new_n544), .B2(G52), .ZN(G171));
  NAND2_X1  g133(.A1(G68), .A2(G543), .ZN(new_n559));
  INV_X1    g134(.A(G56), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n559), .B1(new_n519), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G651), .ZN(new_n562));
  INV_X1    g137(.A(G81), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n562), .B1(new_n563), .B2(new_n556), .ZN(new_n564));
  INV_X1    g139(.A(G43), .ZN(new_n565));
  AOI21_X1  g140(.A(new_n565), .B1(new_n542), .B2(new_n543), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(new_n568));
  XOR2_X1   g143(.A(new_n568), .B(KEYINPUT78), .Z(G153));
  AND3_X1   g144(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G36), .ZN(G176));
  XOR2_X1   g146(.A(KEYINPUT79), .B(KEYINPUT8), .Z(new_n572));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G188));
  NAND2_X1  g150(.A1(G78), .A2(G543), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT80), .ZN(new_n577));
  XOR2_X1   g152(.A(KEYINPUT81), .B(G65), .Z(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n519), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(new_n534), .B2(G91), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n528), .A2(G53), .A3(G543), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(KEYINPUT9), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT9), .ZN(new_n583));
  NAND4_X1  g158(.A1(new_n528), .A2(new_n583), .A3(G53), .A4(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n580), .A2(new_n585), .ZN(G299));
  INV_X1    g161(.A(G171), .ZN(G301));
  NAND2_X1  g162(.A1(new_n530), .A2(G49), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n534), .A2(G87), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n588), .A2(new_n589), .A3(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G61), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n519), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n530), .A2(G48), .B1(new_n594), .B2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n534), .A2(G86), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(G305));
  AND2_X1   g173(.A1(new_n544), .A2(G47), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G651), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  OAI22_X1  g177(.A1(new_n600), .A2(new_n601), .B1(new_n556), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n544), .A2(G54), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n534), .A2(KEYINPUT10), .A3(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  INV_X1    g184(.A(G92), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n556), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n515), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(new_n601), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n607), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n606), .B1(G868), .B2(new_n616), .ZN(G284));
  XNOR2_X1  g192(.A(G284), .B(KEYINPUT82), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  XOR2_X1   g194(.A(G299), .B(KEYINPUT83), .Z(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT84), .ZN(G148));
  NAND2_X1  g200(.A1(new_n616), .A2(new_n623), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G868), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G868), .B2(new_n567), .ZN(G323));
  XNOR2_X1  g203(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g204(.A(new_n475), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(new_n504), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(KEYINPUT12), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2100), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n482), .A2(G123), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT85), .ZN(new_n636));
  INV_X1    g211(.A(new_n470), .ZN(new_n637));
  INV_X1    g212(.A(G135), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  OR2_X1    g214(.A1(G99), .A2(G2105), .ZN(new_n640));
  OAI211_X1 g215(.A(new_n640), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n470), .A2(KEYINPUT85), .A3(G135), .ZN(new_n642));
  AND4_X1   g217(.A1(new_n635), .A2(new_n639), .A3(new_n641), .A4(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2096), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n634), .A2(new_n644), .ZN(G156));
  XOR2_X1   g220(.A(KEYINPUT15), .B(G2435), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2438), .ZN(new_n647));
  XOR2_X1   g222(.A(G2427), .B(G2430), .Z(new_n648));
  OAI21_X1  g223(.A(KEYINPUT14), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT87), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n648), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G2451), .B(G2454), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(G2443), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2446), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G1341), .B(G1348), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n657), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n659), .B1(new_n657), .B2(new_n660), .ZN(new_n662));
  XNOR2_X1  g237(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  OR3_X1    g239(.A1(new_n661), .A2(new_n662), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n664), .B1(new_n661), .B2(new_n662), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n667), .A2(KEYINPUT88), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(KEYINPUT88), .ZN(new_n669));
  AND2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(G401));
  XOR2_X1   g245(.A(G2084), .B(G2090), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT89), .ZN(new_n672));
  XOR2_X1   g247(.A(G2067), .B(G2678), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2072), .B(G2078), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT18), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n675), .B(KEYINPUT17), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n679), .A2(new_n673), .A3(new_n672), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT90), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n672), .B1(new_n674), .B2(new_n678), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n682), .B1(new_n674), .B2(new_n675), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n677), .A2(new_n681), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT91), .B(G2096), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G2100), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n684), .B(new_n686), .ZN(G227));
  XNOR2_X1  g262(.A(G1971), .B(G1976), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT19), .ZN(new_n689));
  XOR2_X1   g264(.A(G1956), .B(G2474), .Z(new_n690));
  XOR2_X1   g265(.A(G1961), .B(G1966), .Z(new_n691));
  NAND2_X1  g266(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT92), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n690), .A2(new_n691), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(new_n692), .ZN(new_n699));
  MUX2_X1   g274(.A(new_n698), .B(new_n699), .S(new_n689), .Z(new_n700));
  NAND2_X1  g275(.A1(new_n696), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1991), .B(G1996), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(G1981), .B(G1986), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT93), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n705), .B(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(G229));
  OR2_X1    g284(.A1(G16), .A2(G21), .ZN(new_n710));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(G286), .B2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G1966), .ZN(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT30), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n715), .A2(G28), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(G28), .ZN(new_n717));
  AND2_X1   g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  AOI22_X1  g293(.A1(new_n712), .A2(new_n713), .B1(new_n714), .B2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT31), .B(G11), .ZN(new_n720));
  NAND2_X1  g295(.A1(G171), .A2(G16), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n721), .B(G1961), .C1(G5), .C2(G16), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n719), .A2(new_n720), .A3(new_n722), .ZN(new_n723));
  OAI211_X1 g298(.A(G1966), .B(new_n710), .C1(G286), .C2(new_n711), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT102), .Z(new_n725));
  INV_X1    g300(.A(KEYINPUT103), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n643), .A2(G29), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n723), .A2(new_n725), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n719), .A2(new_n727), .A3(new_n720), .A4(new_n722), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n724), .B(KEYINPUT102), .ZN(new_n730));
  OAI21_X1  g305(.A(KEYINPUT103), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT28), .ZN(new_n733));
  INV_X1    g308(.A(G26), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(G29), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n734), .A2(G29), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT97), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n482), .A2(new_n737), .A3(G128), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n504), .A2(G2105), .ZN(new_n739));
  INV_X1    g314(.A(G128), .ZN(new_n740));
  OAI21_X1  g315(.A(KEYINPUT97), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n470), .A2(G140), .ZN(new_n742));
  OR2_X1    g317(.A1(G104), .A2(G2105), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n743), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n738), .A2(new_n741), .A3(new_n742), .A4(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(KEYINPUT98), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n742), .A2(new_n744), .ZN(new_n747));
  INV_X1    g322(.A(KEYINPUT98), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n747), .A2(new_n748), .A3(new_n741), .A4(new_n738), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n736), .B1(new_n750), .B2(G29), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n735), .B1(new_n751), .B2(new_n733), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n752), .A2(G2067), .ZN(new_n753));
  NAND3_X1  g328(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT100), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT26), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n482), .A2(G129), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n630), .A2(G105), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n470), .A2(G141), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NOR3_X1   g336(.A1(new_n757), .A2(new_n761), .A3(new_n714), .ZN(new_n762));
  NOR2_X1   g337(.A1(G29), .A2(G32), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT27), .B(G1996), .Z(new_n765));
  OAI21_X1  g340(.A(KEYINPUT101), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT101), .ZN(new_n767));
  INV_X1    g342(.A(new_n765), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n767), .B(new_n768), .C1(new_n762), .C2(new_n763), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n721), .B1(G5), .B2(G16), .ZN(new_n770));
  INV_X1    g345(.A(G1961), .ZN(new_n771));
  AOI22_X1  g346(.A1(new_n766), .A2(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n764), .A2(new_n765), .ZN(new_n773));
  INV_X1    g348(.A(G2067), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n774), .B(new_n735), .C1(new_n751), .C2(new_n733), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n753), .A2(new_n772), .A3(new_n773), .A4(new_n775), .ZN(new_n776));
  NOR2_X1   g351(.A1(G27), .A2(G29), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n777), .B1(G164), .B2(G29), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n778), .A2(G2078), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n714), .A2(G35), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G162), .B2(new_n714), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT104), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT29), .ZN(new_n784));
  AOI22_X1  g359(.A1(new_n784), .A2(G2090), .B1(G2078), .B2(new_n778), .ZN(new_n785));
  OR2_X1    g360(.A1(G29), .A2(G33), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT25), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n470), .A2(G139), .ZN(new_n789));
  AOI22_X1  g364(.A1(new_n504), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n788), .B(new_n789), .C1(new_n469), .C2(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n786), .B1(new_n791), .B2(new_n714), .ZN(new_n792));
  INV_X1    g367(.A(G2072), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n732), .A2(new_n780), .A3(new_n785), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n711), .A2(G4), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(new_n616), .B2(new_n711), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(G1348), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n784), .A2(G2090), .ZN(new_n799));
  NOR3_X1   g374(.A1(new_n795), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n792), .A2(new_n793), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(KEYINPUT99), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n711), .A2(G19), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n567), .B2(new_n711), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G1341), .Z(new_n805));
  NAND3_X1  g380(.A1(new_n711), .A2(KEYINPUT23), .A3(G20), .ZN(new_n806));
  INV_X1    g381(.A(KEYINPUT23), .ZN(new_n807));
  INV_X1    g382(.A(G20), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n807), .B1(new_n808), .B2(G16), .ZN(new_n809));
  INV_X1    g384(.A(G299), .ZN(new_n810));
  OAI211_X1 g385(.A(new_n806), .B(new_n809), .C1(new_n810), .C2(new_n711), .ZN(new_n811));
  INV_X1    g386(.A(G1956), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n800), .A2(new_n802), .A3(new_n805), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n711), .A2(G6), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n597), .B2(new_n711), .ZN(new_n816));
  XOR2_X1   g391(.A(KEYINPUT32), .B(G1981), .Z(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT96), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n816), .B(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n711), .A2(G22), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G303), .B2(G16), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(G1971), .ZN(new_n822));
  NOR2_X1   g397(.A1(G16), .A2(G23), .ZN(new_n823));
  INV_X1    g398(.A(G288), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n823), .B1(new_n824), .B2(G16), .ZN(new_n825));
  XNOR2_X1  g400(.A(KEYINPUT33), .B(G1976), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n819), .A2(new_n822), .A3(new_n827), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT34), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n714), .A2(G25), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n482), .A2(G119), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT94), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n470), .A2(G131), .ZN(new_n833));
  NOR2_X1   g408(.A1(G95), .A2(G2105), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(new_n469), .B2(G107), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n832), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n830), .B1(new_n837), .B2(new_n714), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT35), .B(G1991), .Z(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT95), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n838), .B(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n711), .A2(G24), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n604), .B2(new_n711), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(G1986), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n829), .A2(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n846), .A2(KEYINPUT36), .ZN(new_n847));
  NOR2_X1   g422(.A1(new_n846), .A2(KEYINPUT36), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  OR2_X1    g424(.A1(KEYINPUT24), .A2(G34), .ZN(new_n850));
  NAND2_X1  g425(.A1(KEYINPUT24), .A2(G34), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(new_n714), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(G160), .B2(new_n714), .ZN(new_n853));
  INV_X1    g428(.A(G2084), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n814), .A2(new_n849), .A3(new_n856), .ZN(G311));
  AND3_X1   g432(.A1(new_n800), .A2(new_n805), .A3(new_n813), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n847), .A2(new_n848), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n858), .A2(new_n859), .A3(new_n855), .A4(new_n802), .ZN(G150));
  NAND2_X1  g435(.A1(G80), .A2(G543), .ZN(new_n861));
  INV_X1    g436(.A(G67), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n519), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(G651), .ZN(new_n864));
  INV_X1    g439(.A(G93), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n864), .B1(new_n865), .B2(new_n556), .ZN(new_n866));
  INV_X1    g441(.A(G55), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n542), .B2(new_n543), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(G860), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(KEYINPUT106), .B(KEYINPUT37), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n544), .A2(G43), .ZN(new_n874));
  AOI22_X1  g449(.A1(new_n534), .A2(G81), .B1(new_n561), .B2(G651), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n874), .B(new_n875), .C1(new_n868), .C2(new_n866), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n544), .A2(G55), .ZN(new_n877));
  AOI22_X1  g452(.A1(new_n534), .A2(G93), .B1(new_n863), .B2(G651), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n877), .B(new_n878), .C1(new_n566), .C2(new_n564), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n876), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT38), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n616), .A2(G559), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(KEYINPUT39), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT105), .Z(new_n885));
  OAI21_X1  g460(.A(new_n870), .B1(new_n883), .B2(KEYINPUT39), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n873), .B1(new_n885), .B2(new_n886), .ZN(G145));
  XNOR2_X1  g462(.A(new_n750), .B(new_n632), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n837), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n757), .A2(new_n761), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(new_n791), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n889), .B(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n487), .B(KEYINPUT107), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(G160), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(new_n643), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n482), .A2(G130), .B1(new_n470), .B2(G142), .ZN(new_n896));
  OAI21_X1  g471(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  OAI211_X1 g475(.A(new_n899), .B(new_n900), .C1(G118), .C2(new_n469), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  XOR2_X1   g477(.A(new_n902), .B(new_n509), .Z(new_n903));
  XNOR2_X1  g478(.A(new_n895), .B(new_n903), .ZN(new_n904));
  OR2_X1    g479(.A1(new_n892), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n892), .A2(new_n904), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  XNOR2_X1  g483(.A(new_n908), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g484(.A1(new_n615), .A2(G559), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n880), .B(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n615), .A2(G299), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n616), .A2(new_n810), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n914), .A2(KEYINPUT109), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n912), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT41), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n913), .A2(KEYINPUT41), .A3(new_n912), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OR2_X1    g495(.A1(new_n920), .A2(new_n911), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n914), .A2(KEYINPUT109), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n915), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT42), .ZN(new_n924));
  NAND2_X1  g499(.A1(G303), .A2(new_n824), .ZN(new_n925));
  NAND3_X1  g500(.A1(G288), .A2(new_n523), .A3(new_n535), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n597), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(G305), .A3(new_n926), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n928), .A2(new_n604), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g505(.A(new_n604), .B1(new_n928), .B2(new_n929), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n934));
  NAND4_X1  g509(.A1(new_n915), .A2(new_n934), .A3(new_n921), .A4(new_n922), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n924), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n933), .B1(new_n924), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(G868), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n938), .B1(G868), .B2(new_n869), .ZN(G295));
  OAI21_X1  g514(.A(new_n938), .B1(G868), .B2(new_n869), .ZN(G331));
  NAND3_X1  g515(.A1(new_n876), .A2(new_n879), .A3(G286), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(G286), .B1(new_n876), .B2(new_n879), .ZN(new_n943));
  OAI21_X1  g518(.A(G301), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n880), .A2(G168), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(G171), .A3(new_n941), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n944), .A2(new_n916), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  AOI22_X1  g524(.A1(new_n944), .A2(new_n946), .B1(new_n918), .B2(new_n919), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n933), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n944), .A2(new_n946), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(new_n920), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n953), .A2(new_n948), .A3(new_n932), .A4(new_n947), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n951), .A2(new_n906), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n951), .A2(new_n954), .A3(new_n957), .A4(new_n906), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n956), .A2(KEYINPUT111), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n958), .A2(KEYINPUT111), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT44), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n956), .A2(new_n958), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n961), .A2(new_n964), .ZN(G397));
  INV_X1    g540(.A(G1384), .ZN(new_n966));
  AOI22_X1  g541(.A1(new_n504), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n967));
  OAI22_X1  g542(.A1(new_n967), .A2(new_n469), .B1(new_n490), .B2(new_n489), .ZN(new_n968));
  AND4_X1   g543(.A1(new_n463), .A2(new_n465), .A3(new_n501), .A4(new_n506), .ZN(new_n969));
  AOI22_X1  g544(.A1(new_n969), .A2(new_n497), .B1(new_n502), .B2(new_n499), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n966), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n971), .B(KEYINPUT112), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n471), .A2(new_n480), .A3(G40), .ZN(new_n975));
  NOR2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  NOR3_X1   g552(.A1(new_n977), .A2(G1986), .A3(G290), .ZN(new_n978));
  XOR2_X1   g553(.A(new_n978), .B(KEYINPUT48), .Z(new_n979));
  XNOR2_X1  g554(.A(new_n750), .B(G2067), .ZN(new_n980));
  INV_X1    g555(.A(G1996), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n890), .B(new_n981), .ZN(new_n982));
  OR2_X1    g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  XOR2_X1   g558(.A(new_n837), .B(new_n840), .Z(new_n984));
  OAI21_X1  g559(.A(new_n976), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n979), .A2(new_n985), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n750), .A2(G2067), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n983), .A2(new_n976), .ZN(new_n988));
  INV_X1    g563(.A(new_n837), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(new_n840), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n987), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT126), .ZN(new_n992));
  OR2_X1    g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n991), .A2(new_n992), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n976), .A3(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT46), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(new_n977), .B2(G1996), .ZN(new_n997));
  INV_X1    g572(.A(new_n890), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n976), .B1(new_n998), .B2(new_n980), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n976), .A2(KEYINPUT46), .A3(new_n981), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  XNOR2_X1  g576(.A(new_n1001), .B(KEYINPUT47), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n986), .A2(new_n995), .A3(new_n1002), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n971), .A2(new_n975), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT114), .B(G8), .Z(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n824), .A2(G1976), .ZN(new_n1008));
  AOI21_X1  g583(.A(KEYINPUT52), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n824), .B2(G1976), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1007), .B(new_n1011), .C1(KEYINPUT52), .C2(new_n1008), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT117), .B(G86), .Z(new_n1015));
  OAI21_X1  g590(.A(new_n595), .B1(new_n556), .B2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(G1981), .ZN(new_n1017));
  XOR2_X1   g592(.A(KEYINPUT116), .B(G1981), .Z(new_n1018));
  NAND3_X1  g593(.A1(new_n595), .A2(new_n596), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(KEYINPUT49), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT49), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1013), .A2(new_n1014), .B1(new_n1023), .B2(new_n1007), .ZN(new_n1024));
  NAND2_X1  g599(.A1(G303), .A2(G8), .ZN(new_n1025));
  XOR2_X1   g600(.A(new_n1025), .B(KEYINPUT55), .Z(new_n1026));
  INV_X1    g601(.A(KEYINPUT50), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n971), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1384), .B1(new_n495), .B2(new_n508), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT50), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n975), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(G2090), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n971), .A2(new_n973), .ZN(new_n1034));
  INV_X1    g609(.A(new_n975), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1029), .A2(KEYINPUT45), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(G1971), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1033), .A2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1024), .A2(G8), .A3(new_n1026), .A4(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1022), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1042), .A2(new_n1007), .A3(new_n1020), .ZN(new_n1043));
  INV_X1    g618(.A(G1976), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1043), .A2(new_n1044), .A3(new_n824), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n1019), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1046), .A2(KEYINPUT119), .ZN(new_n1047));
  XNOR2_X1  g622(.A(new_n1007), .B(KEYINPUT118), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1046), .A2(KEYINPUT119), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1006), .B1(new_n1033), .B2(new_n1039), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1051), .A2(new_n1026), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1026), .A2(new_n1040), .A3(G8), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1052), .A2(new_n1024), .A3(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT120), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1034), .A2(KEYINPUT120), .A3(new_n1035), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1036), .A3(new_n1058), .ZN(new_n1059));
  AOI22_X1  g634(.A1(new_n1059), .A2(new_n713), .B1(new_n854), .B2(new_n1031), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1060), .A2(G286), .A3(new_n1006), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT63), .B1(new_n1054), .B2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1026), .B1(G8), .B2(new_n1040), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  AND4_X1   g640(.A1(new_n1053), .A2(new_n1061), .A3(new_n1065), .A4(new_n1024), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n1041), .B(new_n1050), .C1(new_n1062), .C2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(G168), .A2(new_n1006), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G8), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1069), .B1(new_n1060), .B2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1071), .A2(KEYINPUT51), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1068), .A2(KEYINPUT51), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1073), .B1(new_n1060), .B2(new_n1006), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1060), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1068), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1037), .B2(G2078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT50), .B1(new_n509), .B2(new_n966), .ZN(new_n1080));
  AOI211_X1 g655(.A(new_n1027), .B(G1384), .C1(new_n495), .C2(new_n508), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1035), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT123), .B(G1961), .Z(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G2078), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(KEYINPUT53), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n1079), .B(new_n1084), .C1(new_n1059), .C2(new_n1086), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1087), .A2(KEYINPUT62), .A3(G171), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1075), .A2(new_n1077), .A3(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1087), .A2(G171), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1090), .A2(KEYINPUT62), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT122), .B(G2072), .ZN(new_n1092));
  XNOR2_X1  g667(.A(new_n1092), .B(KEYINPUT56), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n579), .A2(G651), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n534), .A2(G91), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(KEYINPUT121), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n1098));
  NAND3_X1  g673(.A1(G299), .A2(new_n1097), .A3(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n580), .B(new_n585), .C1(KEYINPUT121), .C2(KEYINPUT57), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI211_X1 g676(.A(new_n1094), .B(new_n1101), .C1(new_n1031), .C2(G1956), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1082), .A2(new_n812), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1101), .B1(new_n1103), .B2(new_n1094), .ZN(new_n1104));
  INV_X1    g679(.A(G1348), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1082), .A2(new_n1105), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n971), .A2(new_n975), .A3(G2067), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n615), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1102), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  AOI211_X1 g685(.A(new_n616), .B(new_n1107), .C1(new_n1082), .C2(new_n1105), .ZN(new_n1111));
  OAI21_X1  g686(.A(KEYINPUT60), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1034), .A2(new_n981), .A3(new_n1036), .A4(new_n1035), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT58), .B(G1341), .Z(new_n1114));
  OAI21_X1  g689(.A(new_n1114), .B1(new_n971), .B2(new_n975), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT59), .B1(new_n1116), .B2(new_n567), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n1118));
  INV_X1    g693(.A(new_n567), .ZN(new_n1119));
  AOI211_X1 g694(.A(new_n1118), .B(new_n1119), .C1(new_n1113), .C2(new_n1115), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1117), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1106), .A2(new_n1122), .A3(new_n616), .A4(new_n1108), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1112), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT61), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1102), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(new_n1126), .B2(new_n1104), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1094), .B1(new_n1031), .B2(G1956), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1101), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(KEYINPUT61), .A3(new_n1102), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1127), .A2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1110), .B1(new_n1124), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1035), .B1(KEYINPUT124), .B2(new_n1085), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(KEYINPUT124), .B2(new_n1085), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1135), .A2(new_n974), .A3(KEYINPUT53), .A4(new_n1036), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1136), .A2(new_n1079), .A3(new_n1084), .ZN(new_n1137));
  XOR2_X1   g712(.A(G171), .B(KEYINPUT54), .Z(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1087), .B2(new_n1139), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1091), .B1(new_n1133), .B2(new_n1141), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1072), .A2(new_n1074), .B1(new_n1076), .B2(new_n1068), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1089), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(new_n1054), .B(KEYINPUT125), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1067), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n604), .B(G1986), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n985), .B1(new_n977), .B2(new_n1147), .ZN(new_n1148));
  XOR2_X1   g723(.A(new_n1148), .B(KEYINPUT113), .Z(new_n1149));
  OAI21_X1  g724(.A(new_n1003), .B1(new_n1146), .B2(new_n1149), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g725(.A1(G227), .A2(new_n459), .ZN(new_n1152));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n1153));
  NOR2_X1   g727(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g728(.A(new_n1154), .B1(new_n668), .B2(new_n669), .ZN(new_n1155));
  AOI22_X1  g729(.A1(new_n956), .A2(new_n958), .B1(new_n1153), .B2(new_n1152), .ZN(new_n1156));
  AND4_X1   g730(.A1(new_n708), .A2(new_n1155), .A3(new_n908), .A4(new_n1156), .ZN(G308));
  NAND4_X1  g731(.A1(new_n708), .A2(new_n1155), .A3(new_n908), .A4(new_n1156), .ZN(G225));
endmodule


