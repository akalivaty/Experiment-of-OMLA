//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(KEYINPUT16), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND3_X1  g002(.A1(new_n187), .A2(new_n188), .A3(G125), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G125), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n189), .B1(new_n193), .B2(new_n187), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI211_X1 g010(.A(G146), .B(new_n189), .C1(new_n193), .C2(new_n187), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(G128), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G119), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT24), .B(G110), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT23), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n201), .A2(KEYINPUT23), .A3(G119), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n200), .A3(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n205), .B1(G110), .B2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n198), .A2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G110), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n207), .A2(new_n208), .A3(new_n212), .A4(new_n200), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT71), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n203), .A2(new_n204), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n213), .B2(new_n214), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT72), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n197), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(G125), .B(G140), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(KEYINPUT16), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n222), .A2(KEYINPUT72), .A3(G146), .A4(new_n189), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n221), .A2(new_n195), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n220), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n211), .B1(new_n218), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT22), .B(G137), .ZN(new_n227));
  INV_X1    g041(.A(G953), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(G221), .A3(G234), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n227), .B(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n226), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G902), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n211), .B(new_n230), .C1(new_n218), .C2(new_n225), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n232), .A2(KEYINPUT25), .A3(new_n233), .A4(new_n234), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G217), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n240), .B1(G234), .B2(new_n233), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n232), .A2(new_n234), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n241), .A2(G902), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n239), .A2(new_n241), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n247));
  INV_X1    g061(.A(G237), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(new_n228), .A3(G210), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n249), .B(KEYINPUT27), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G101), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT68), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT11), .ZN(new_n254));
  INV_X1    g068(.A(G134), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n254), .B1(new_n255), .B2(G137), .ZN(new_n256));
  INV_X1    g070(.A(G137), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(KEYINPUT11), .A3(G134), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(G137), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n256), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G131), .ZN(new_n261));
  INV_X1    g075(.A(G131), .ZN(new_n262));
  NAND4_X1  g076(.A1(new_n256), .A2(new_n258), .A3(new_n262), .A4(new_n259), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(KEYINPUT0), .A2(G128), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(G143), .B(G146), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n268), .B1(KEYINPUT0), .B2(G128), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n266), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT0), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT65), .B1(new_n271), .B2(new_n201), .ZN(new_n272));
  INV_X1    g086(.A(G143), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n273), .A2(G146), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n195), .A2(G143), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n272), .B(new_n265), .C1(new_n274), .C2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n253), .B1(new_n264), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G113), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT2), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT2), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G113), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT67), .B1(new_n199), .B2(G116), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT67), .ZN(new_n285));
  INV_X1    g099(.A(G116), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(new_n286), .A3(G119), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n286), .A2(G119), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n283), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(KEYINPUT1), .B1(new_n273), .B2(G146), .ZN(new_n293));
  OAI211_X1 g107(.A(G128), .B(new_n293), .C1(new_n274), .C2(new_n275), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n255), .A2(G137), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n257), .A2(G134), .ZN(new_n296));
  OAI21_X1  g110(.A(G131), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n195), .A2(G143), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n273), .A2(G146), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n298), .B(new_n299), .C1(KEYINPUT1), .C2(new_n201), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n294), .A2(new_n263), .A3(new_n297), .A4(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n288), .A2(new_n290), .A3(new_n283), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n292), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(new_n277), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n261), .A2(new_n263), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(KEYINPUT68), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n278), .A2(new_n303), .A3(new_n306), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n288), .A2(new_n290), .A3(new_n283), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n308), .A2(new_n291), .ZN(new_n309));
  INV_X1    g123(.A(new_n301), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT66), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n277), .A2(new_n311), .B1(new_n263), .B2(new_n261), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n270), .A2(new_n276), .A3(KEYINPUT66), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n310), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n307), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT28), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n304), .A2(new_n305), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n303), .A2(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n318), .A2(KEYINPUT28), .ZN(new_n319));
  INV_X1    g133(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n252), .B1(new_n316), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT31), .ZN(new_n322));
  INV_X1    g136(.A(new_n309), .ZN(new_n323));
  XNOR2_X1  g137(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n323), .B1(new_n314), .B2(new_n324), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n301), .A2(KEYINPUT30), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n278), .A2(new_n306), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT69), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n278), .A2(new_n306), .A3(KEYINPUT69), .A4(new_n326), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n325), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n307), .A2(new_n252), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n322), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n329), .A2(new_n330), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n312), .A2(new_n313), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(new_n301), .ZN(new_n336));
  INV_X1    g150(.A(new_n324), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n309), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n332), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(KEYINPUT31), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n321), .B1(new_n333), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(G472), .A2(G902), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n247), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n321), .ZN(new_n346));
  AOI21_X1  g160(.A(KEYINPUT31), .B1(new_n339), .B2(new_n340), .ZN(new_n347));
  AOI211_X1 g161(.A(new_n322), .B(new_n332), .C1(new_n334), .C2(new_n338), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n346), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(KEYINPUT70), .A3(new_n343), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n345), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(G472), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n316), .A2(new_n320), .A3(new_n252), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT29), .ZN(new_n355));
  INV_X1    g169(.A(new_n307), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n356), .B1(new_n334), .B2(new_n338), .ZN(new_n357));
  OAI211_X1 g171(.A(new_n354), .B(new_n355), .C1(new_n357), .C2(new_n252), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n278), .A2(new_n301), .A3(new_n306), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n323), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n307), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n319), .B1(new_n361), .B2(KEYINPUT28), .ZN(new_n362));
  INV_X1    g176(.A(new_n252), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(new_n355), .ZN(new_n364));
  AOI21_X1  g178(.A(G902), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n353), .B1(new_n358), .B2(new_n365), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n342), .A2(new_n344), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n366), .B1(new_n367), .B2(KEYINPUT32), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n246), .B1(new_n352), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(G113), .B(G122), .ZN(new_n370));
  INV_X1    g184(.A(G104), .ZN(new_n371));
  XNOR2_X1  g185(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n248), .A2(new_n228), .A3(G214), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT85), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n374), .B1(KEYINPUT84), .B2(G143), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n273), .A2(KEYINPUT85), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AND3_X1   g191(.A1(new_n248), .A2(new_n228), .A3(G214), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT84), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT85), .B1(new_n379), .B2(new_n273), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  OAI211_X1 g195(.A(KEYINPUT18), .B(G131), .C1(new_n377), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n193), .A2(G146), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(new_n224), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n374), .A2(G143), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n378), .B1(new_n380), .B2(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n386), .B1(new_n380), .B2(new_n378), .ZN(new_n387));
  AND2_X1   g201(.A1(KEYINPUT18), .A2(G131), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n382), .B(new_n384), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(new_n386), .B(new_n262), .C1(new_n380), .C2(new_n378), .ZN(new_n390));
  OAI21_X1  g204(.A(G131), .B1(new_n377), .B2(new_n381), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT17), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n390), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n197), .B(new_n196), .C1(new_n391), .C2(new_n392), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n372), .B(new_n389), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n390), .A2(new_n391), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT86), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n398), .B(KEYINPUT19), .C1(new_n193), .C2(KEYINPUT87), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT87), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT86), .B1(new_n221), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT19), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n402), .B1(new_n221), .B2(KEYINPUT86), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n399), .B(new_n195), .C1(new_n401), .C2(new_n403), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n397), .A2(new_n220), .A3(new_n223), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n372), .B1(new_n405), .B2(new_n389), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n396), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(G475), .A2(G902), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT20), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT88), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n412), .B1(new_n396), .B2(new_n406), .ZN(new_n413));
  AND2_X1   g227(.A1(new_n405), .A2(new_n389), .ZN(new_n414));
  OAI211_X1 g228(.A(KEYINPUT88), .B(new_n395), .C1(new_n414), .C2(new_n372), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n415), .A3(new_n408), .ZN(new_n416));
  XNOR2_X1  g230(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n411), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  XNOR2_X1  g233(.A(G128), .B(G143), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT13), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n201), .A2(KEYINPUT13), .A3(G143), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(new_n255), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n255), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT91), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n421), .A2(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n286), .A2(G122), .ZN(new_n427));
  INV_X1    g241(.A(G122), .ZN(new_n428));
  OAI21_X1  g242(.A(KEYINPUT90), .B1(new_n428), .B2(G116), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT90), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n286), .A3(G122), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n427), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(G107), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n432), .A2(new_n433), .ZN(new_n436));
  OAI221_X1 g250(.A(new_n426), .B1(new_n425), .B2(new_n424), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT9), .B(G234), .ZN(new_n438));
  NOR3_X1   g252(.A1(new_n438), .A2(new_n240), .A3(G953), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n429), .A2(new_n431), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n427), .B1(new_n440), .B2(KEYINPUT14), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT14), .ZN(new_n442));
  AND2_X1   g256(.A1(new_n429), .A2(new_n431), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n441), .A2(KEYINPUT93), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT93), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n442), .B1(new_n429), .B2(new_n431), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n445), .B1(new_n446), .B2(new_n427), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n433), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n420), .A2(new_n255), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n424), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT92), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n432), .A2(new_n451), .A3(new_n433), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n451), .B1(new_n432), .B2(new_n433), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n450), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n437), .B(new_n439), .C1(new_n448), .C2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n427), .ZN(new_n458));
  OAI211_X1 g272(.A(KEYINPUT93), .B(new_n458), .C1(new_n443), .C2(new_n442), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n443), .A2(new_n442), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n459), .A2(new_n447), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(G107), .ZN(new_n462));
  INV_X1    g276(.A(new_n454), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n463), .A2(new_n452), .B1(new_n424), .B2(new_n449), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n439), .B1(new_n465), .B2(new_n437), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n233), .B1(new_n457), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G478), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n468), .A2(KEYINPUT15), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n437), .B1(new_n448), .B2(new_n455), .ZN(new_n471));
  INV_X1    g285(.A(new_n439), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(G902), .B1(new_n473), .B2(new_n456), .ZN(new_n474));
  INV_X1    g288(.A(new_n469), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g290(.A1(new_n228), .A2(G952), .ZN(new_n477));
  INV_X1    g291(.A(G234), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n477), .B1(new_n478), .B2(new_n248), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(G902), .B(G953), .C1(new_n478), .C2(new_n248), .ZN(new_n481));
  XNOR2_X1  g295(.A(new_n481), .B(KEYINPUT94), .ZN(new_n482));
  XNOR2_X1  g296(.A(KEYINPUT21), .B(G898), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n470), .A2(new_n476), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G475), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n389), .B1(new_n393), .B2(new_n394), .ZN(new_n488));
  INV_X1    g302(.A(new_n372), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT89), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n492), .A2(G902), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(new_n491), .A3(new_n395), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n487), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n419), .A2(new_n486), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G214), .B1(G237), .B2(G902), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n288), .A2(KEYINPUT5), .A3(new_n290), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT5), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n279), .B1(new_n289), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(KEYINPUT3), .B1(new_n371), .B2(G107), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT3), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n504), .A2(new_n433), .A3(G104), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n433), .A2(G104), .ZN(new_n507));
  AND2_X1   g321(.A1(KEYINPUT76), .A2(G101), .ZN(new_n508));
  NOR2_X1   g322(.A1(KEYINPUT76), .A2(G101), .ZN(new_n509));
  NOR3_X1   g323(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n371), .A2(G107), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n433), .A2(G104), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g327(.A1(new_n506), .A2(new_n510), .B1(G101), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n502), .A2(new_n514), .A3(new_n302), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n503), .A2(new_n505), .A3(new_n511), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT4), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n517), .A3(G101), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n518), .B1(new_n308), .B2(new_n291), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(G101), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n508), .A2(new_n509), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n521), .A2(new_n511), .A3(new_n503), .A4(new_n505), .ZN(new_n522));
  AND3_X1   g336(.A1(new_n520), .A2(KEYINPUT4), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n515), .B1(new_n519), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g338(.A(G110), .B(G122), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n515), .B(new_n525), .C1(new_n519), .C2(new_n523), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n527), .A2(KEYINPUT6), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n277), .A2(G125), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT80), .B(G224), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n228), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n294), .A2(new_n300), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(new_n191), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n530), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n532), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n191), .B1(new_n270), .B2(new_n276), .ZN(new_n537));
  AOI21_X1  g351(.A(G125), .B1(new_n294), .B2(new_n300), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT6), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n524), .A2(new_n541), .A3(new_n526), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n529), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n233), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT7), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n532), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n547), .B1(new_n530), .B2(new_n534), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n540), .B2(new_n547), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n525), .B(KEYINPUT8), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n502), .A2(new_n514), .A3(new_n302), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n514), .B1(new_n502), .B2(new_n302), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT81), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n532), .B1(new_n530), .B2(new_n534), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n537), .A2(new_n538), .A3(new_n536), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n547), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n548), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n559), .A2(KEYINPUT81), .A3(new_n553), .A4(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n556), .A2(new_n528), .A3(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(G210), .B1(G237), .B2(G902), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n545), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(KEYINPUT82), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n528), .ZN(new_n566));
  AOI21_X1  g380(.A(KEYINPUT81), .B1(new_n549), .B2(new_n553), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n565), .B1(new_n568), .B2(new_n544), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n498), .B1(new_n564), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G469), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n520), .A2(KEYINPUT4), .A3(new_n522), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n304), .A2(new_n572), .A3(new_n518), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT10), .ZN(new_n574));
  INV_X1    g388(.A(new_n533), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(new_n514), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n513), .A2(G101), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n522), .A2(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n578), .A2(new_n533), .A3(KEYINPUT10), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n264), .B(new_n573), .C1(new_n576), .C2(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT77), .B1(new_n261), .B2(new_n263), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n578), .A2(new_n533), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n522), .A2(new_n577), .B1(new_n294), .B2(new_n300), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT12), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT12), .ZN(new_n586));
  OAI211_X1 g400(.A(new_n586), .B(new_n581), .C1(new_n582), .C2(new_n583), .ZN(new_n587));
  XNOR2_X1  g401(.A(G110), .B(G140), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n228), .A2(G227), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n588), .B(new_n589), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(new_n592));
  AND4_X1   g406(.A1(new_n580), .A2(new_n585), .A3(new_n587), .A4(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n573), .B1(new_n576), .B2(new_n579), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n305), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n592), .B1(new_n595), .B2(new_n580), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n571), .B(new_n233), .C1(new_n593), .C2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n585), .A2(new_n580), .A3(new_n587), .ZN(new_n598));
  INV_X1    g412(.A(new_n592), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n580), .A2(KEYINPUT78), .A3(new_n592), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n595), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT78), .B1(new_n580), .B2(new_n592), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n600), .B(G469), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n571), .A2(new_n233), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n597), .A2(new_n604), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT79), .ZN(new_n608));
  OAI21_X1  g422(.A(G221), .B1(new_n438), .B2(G902), .ZN(new_n609));
  XOR2_X1   g423(.A(new_n609), .B(KEYINPUT73), .Z(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n607), .A2(new_n608), .A3(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n608), .B1(new_n607), .B2(new_n611), .ZN(new_n614));
  OAI211_X1 g428(.A(new_n496), .B(new_n570), .C1(new_n613), .C2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n369), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g431(.A(new_n617), .B(new_n521), .Z(G3));
  OAI21_X1  g432(.A(G472), .B1(new_n342), .B2(G902), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n345), .A2(new_n619), .A3(new_n350), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n607), .A2(new_n611), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n621), .A2(KEYINPUT79), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n246), .B1(new_n622), .B2(new_n612), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n563), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n625), .B1(new_n568), .B2(new_n544), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n564), .A2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n485), .A3(new_n497), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n468), .A2(new_n233), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n474), .B2(new_n468), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT33), .B1(new_n457), .B2(new_n466), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT33), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n473), .A2(new_n632), .A3(new_n456), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n631), .A2(G478), .A3(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT95), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n630), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n635), .B1(new_n630), .B2(new_n634), .ZN(new_n637));
  OAI22_X1  g451(.A1(new_n636), .A2(new_n637), .B1(new_n419), .B2(new_n495), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n624), .A2(new_n628), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT34), .B(G104), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  AND2_X1   g455(.A1(new_n470), .A2(new_n476), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(new_n495), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n416), .A2(new_n418), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n413), .A2(new_n415), .A3(new_n408), .A4(new_n417), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n644), .A2(KEYINPUT96), .A3(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(KEYINPUT96), .B1(new_n644), .B2(new_n645), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n643), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n648), .A2(new_n628), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n649), .A2(new_n620), .A3(new_n623), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT35), .B(G107), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  OAI21_X1  g466(.A(new_n570), .B1(new_n613), .B2(new_n614), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n345), .A2(new_n619), .A3(new_n350), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n239), .A2(new_n241), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n231), .A2(KEYINPUT36), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n226), .B(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n244), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n496), .A2(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n653), .A2(new_n654), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT37), .B(G110), .ZN(new_n662));
  XOR2_X1   g476(.A(new_n662), .B(KEYINPUT97), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n661), .B(new_n663), .ZN(G12));
  NAND2_X1  g478(.A1(new_n352), .A2(new_n368), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n563), .B1(new_n545), .B2(new_n562), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n568), .A2(new_n544), .A3(new_n625), .ZN(new_n667));
  OAI211_X1 g481(.A(new_n497), .B(new_n659), .C1(new_n666), .C2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n612), .B2(new_n622), .ZN(new_n669));
  INV_X1    g483(.A(G900), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n480), .B1(new_n482), .B2(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  OAI211_X1 g486(.A(new_n643), .B(new_n672), .C1(new_n646), .C2(new_n647), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n665), .A2(new_n669), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  NAND2_X1  g490(.A1(new_n622), .A2(new_n612), .ZN(new_n677));
  XOR2_X1   g491(.A(new_n671), .B(KEYINPUT39), .Z(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n677), .A2(new_n678), .A3(new_n680), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT38), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n564), .A2(new_n569), .A3(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n685), .B1(new_n564), .B2(new_n569), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n470), .A2(new_n476), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n690), .B(new_n497), .C1(new_n419), .C2(new_n495), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n689), .A2(new_n659), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n361), .ZN(new_n693));
  AOI21_X1  g507(.A(G902), .B1(new_n693), .B2(new_n363), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n694), .B1(new_n357), .B2(new_n363), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(G472), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT98), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n349), .A2(KEYINPUT32), .A3(new_n343), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n695), .A2(KEYINPUT98), .A3(G472), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n702), .A2(KEYINPUT99), .A3(new_n352), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT99), .B1(new_n702), .B2(new_n352), .ZN(new_n705));
  OAI211_X1 g519(.A(new_n684), .B(new_n692), .C1(new_n704), .C2(new_n705), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT101), .B(G143), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G45));
  NOR2_X1   g522(.A1(new_n638), .A2(new_n671), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n665), .A2(new_n669), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(KEYINPUT102), .B(G146), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G48));
  INV_X1    g526(.A(new_n593), .ZN(new_n713));
  INV_X1    g527(.A(new_n596), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n571), .B1(new_n715), .B2(new_n233), .ZN(new_n716));
  INV_X1    g530(.A(new_n597), .ZN(new_n717));
  INV_X1    g531(.A(new_n609), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n716), .A2(new_n717), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n628), .A2(new_n638), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n369), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT41), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G113), .ZN(G15));
  NAND4_X1  g537(.A1(new_n665), .A2(new_n649), .A3(new_n245), .A4(new_n719), .ZN(new_n724));
  XOR2_X1   g538(.A(KEYINPUT103), .B(G116), .Z(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(G18));
  INV_X1    g540(.A(new_n660), .ZN(new_n727));
  AND3_X1   g541(.A1(new_n719), .A2(new_n497), .A3(new_n627), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n665), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  INV_X1    g544(.A(new_n627), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n731), .A2(new_n691), .A3(new_n484), .ZN(new_n732));
  OAI22_X1  g546(.A1(new_n347), .A2(new_n348), .B1(new_n252), .B2(new_n362), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n343), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n619), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n732), .A2(new_n735), .A3(new_n245), .A4(new_n719), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  AND3_X1   g551(.A1(new_n619), .A2(new_n734), .A3(new_n659), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n709), .A2(new_n728), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  NAND3_X1  g554(.A1(new_n564), .A2(new_n569), .A3(new_n497), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n607), .A2(new_n609), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n665), .A2(new_n245), .A3(new_n709), .A4(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT42), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n709), .A2(new_n743), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n351), .B1(new_n342), .B2(new_n344), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n358), .A2(new_n365), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(G472), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n747), .A2(new_n699), .A3(new_n749), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n750), .A2(KEYINPUT42), .A3(new_n245), .ZN(new_n751));
  AOI22_X1  g565(.A1(new_n744), .A2(new_n745), .B1(new_n746), .B2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(KEYINPUT104), .B(G131), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G33));
  NAND3_X1  g568(.A1(new_n665), .A2(new_n245), .A3(new_n743), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n673), .A2(KEYINPUT105), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n644), .A2(new_n645), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT96), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n644), .A2(KEYINPUT96), .A3(new_n645), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT105), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n761), .A2(new_n762), .A3(new_n643), .A4(new_n672), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n756), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n755), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n255), .ZN(G36));
  OAI21_X1  g580(.A(new_n600), .B1(new_n602), .B2(new_n603), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT45), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n571), .B1(new_n767), .B2(new_n768), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n605), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  OR3_X1    g585(.A1(new_n771), .A2(KEYINPUT106), .A3(KEYINPUT46), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT106), .B1(new_n771), .B2(KEYINPUT46), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n717), .B1(new_n771), .B2(KEYINPUT46), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n772), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n775), .A2(new_n609), .A3(new_n678), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n741), .B(KEYINPUT107), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n419), .A2(new_n495), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n779), .B1(new_n636), .B2(new_n637), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT43), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT43), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n779), .B(new_n782), .C1(new_n636), .C2(new_n637), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n781), .A2(new_n654), .A3(new_n659), .A4(new_n783), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n784), .A2(KEYINPUT44), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n784), .A2(KEYINPUT44), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n776), .B(new_n778), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  INV_X1    g602(.A(new_n638), .ZN(new_n789));
  INV_X1    g603(.A(new_n741), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n789), .A2(new_n246), .A3(new_n672), .A4(new_n790), .ZN(new_n791));
  OR3_X1    g605(.A1(new_n791), .A2(KEYINPUT109), .A3(new_n665), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT109), .B1(new_n791), .B2(new_n665), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n775), .A2(new_n609), .ZN(new_n795));
  XNOR2_X1  g609(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n796));
  OR2_X1    g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT108), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n795), .B1(new_n798), .B2(KEYINPUT47), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n794), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  XOR2_X1   g614(.A(KEYINPUT110), .B(G140), .Z(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(G42));
  OAI21_X1  g616(.A(new_n245), .B1(new_n613), .B2(new_n614), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n642), .A2(new_n419), .A3(new_n495), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n485), .A3(new_n570), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n803), .A2(new_n805), .A3(new_n654), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT111), .B1(new_n806), .B2(new_n661), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n803), .A2(new_n654), .A3(new_n638), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n570), .A2(new_n485), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n808), .A2(new_n809), .B1(new_n369), .B2(new_n616), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n620), .A2(new_n727), .A3(new_n677), .A4(new_n570), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n620), .A2(new_n623), .A3(new_n809), .A4(new_n804), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n807), .A2(new_n810), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n709), .A2(new_n738), .A3(new_n743), .ZN(new_n816));
  INV_X1    g630(.A(new_n665), .ZN(new_n817));
  AOI22_X1  g631(.A1(new_n239), .A2(new_n241), .B1(new_n244), .B2(new_n657), .ZN(new_n818));
  NOR4_X1   g632(.A1(new_n818), .A2(new_n495), .A3(new_n690), .A4(new_n671), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n677), .A2(new_n761), .A3(new_n790), .A4(new_n819), .ZN(new_n820));
  OAI221_X1 g634(.A(new_n816), .B1(new_n817), .B2(new_n820), .C1(new_n755), .C2(new_n764), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n721), .A2(new_n724), .A3(new_n729), .A4(new_n736), .ZN(new_n822));
  NOR4_X1   g636(.A1(new_n815), .A2(new_n821), .A3(new_n822), .A4(new_n752), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n818), .A2(new_n607), .A3(new_n609), .A4(new_n672), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n731), .A2(new_n691), .A3(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n345), .A2(new_n350), .A3(new_n351), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n825), .B1(new_n826), .B2(new_n701), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n675), .A2(new_n710), .A3(new_n739), .A4(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n828), .B(new_n829), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT53), .B1(new_n823), .B2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n807), .A2(new_n810), .A3(new_n814), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n822), .A2(new_n752), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n816), .B1(new_n817), .B2(new_n820), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n765), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n828), .B(KEYINPUT52), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT54), .B1(new_n831), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n838), .B1(new_n836), .B2(new_n837), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(new_n815), .B2(new_n821), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n813), .B1(new_n811), .B2(new_n812), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n620), .A2(new_n623), .A3(new_n789), .A4(new_n809), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n617), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n847), .A2(new_n835), .A3(KEYINPUT112), .A4(new_n814), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n822), .A2(new_n752), .A3(new_n838), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n843), .A2(new_n830), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n841), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n840), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n704), .A2(new_n705), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n790), .A2(new_n719), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n855), .A2(new_n245), .A3(new_n480), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n636), .A2(new_n637), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n857), .A2(new_n779), .A3(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n735), .A2(new_n245), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n860), .A2(new_n719), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n781), .A2(new_n480), .A3(new_n783), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n687), .A2(new_n688), .A3(new_n497), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT50), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n861), .A2(KEYINPUT50), .A3(new_n862), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n859), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n862), .A2(new_n860), .A3(new_n778), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n797), .A2(new_n799), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n716), .A2(new_n717), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n610), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n870), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n862), .A2(new_n738), .A3(new_n855), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT113), .Z(new_n877));
  NAND4_X1  g691(.A1(new_n869), .A2(new_n875), .A3(KEYINPUT51), .A4(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT51), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n859), .A2(new_n877), .A3(new_n868), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n879), .B1(new_n880), .B2(new_n874), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n862), .A2(new_n728), .A3(new_n860), .ZN(new_n882));
  XOR2_X1   g696(.A(new_n882), .B(KEYINPUT114), .Z(new_n883));
  NAND2_X1  g697(.A1(new_n857), .A2(new_n789), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n246), .B1(new_n368), .B2(new_n747), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n862), .A2(new_n885), .A3(new_n855), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT48), .ZN(new_n887));
  AND4_X1   g701(.A1(new_n477), .A2(new_n883), .A3(new_n884), .A4(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n878), .A2(new_n881), .A3(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n853), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  INV_X1    g705(.A(new_n854), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n872), .B(KEYINPUT49), .ZN(new_n893));
  INV_X1    g707(.A(new_n780), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n246), .A2(new_n610), .A3(new_n498), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n893), .A2(new_n689), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  OAI22_X1  g710(.A1(new_n890), .A2(new_n891), .B1(new_n892), .B2(new_n896), .ZN(G75));
  NAND2_X1  g711(.A1(new_n841), .A2(new_n850), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT116), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n898), .A2(new_n899), .A3(G902), .A4(new_n565), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n529), .A2(new_n542), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT115), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT55), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(new_n540), .Z(new_n904));
  INV_X1    g718(.A(KEYINPUT56), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n900), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n233), .B1(new_n841), .B2(new_n850), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n899), .B1(new_n908), .B2(new_n565), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n228), .A2(G952), .ZN(new_n911));
  INV_X1    g725(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(KEYINPUT56), .B1(new_n908), .B2(G210), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n912), .B1(new_n913), .B2(new_n904), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n910), .A2(new_n914), .ZN(G51));
  NAND2_X1  g729(.A1(new_n769), .A2(new_n770), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  AND4_X1   g731(.A1(KEYINPUT117), .A2(new_n898), .A3(G902), .A4(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT117), .B1(new_n908), .B2(new_n917), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n605), .B(KEYINPUT57), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n841), .A2(new_n851), .A3(new_n850), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n851), .B1(new_n841), .B2(new_n850), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n715), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n911), .B1(new_n920), .B2(new_n925), .ZN(G54));
  NAND2_X1  g740(.A1(new_n413), .A2(new_n415), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  AND2_X1   g742(.A1(KEYINPUT58), .A2(G475), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n908), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n928), .B1(new_n908), .B2(new_n929), .ZN(new_n931));
  NOR3_X1   g745(.A1(new_n930), .A2(new_n931), .A3(new_n911), .ZN(G60));
  NAND2_X1  g746(.A1(new_n631), .A2(new_n633), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n629), .B(KEYINPUT59), .Z(new_n934));
  AOI21_X1  g748(.A(new_n933), .B1(new_n853), .B2(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n933), .A2(new_n934), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n936), .B1(new_n922), .B2(new_n923), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n912), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n935), .A2(new_n938), .ZN(G63));
  NAND2_X1  g753(.A1(G217), .A2(G902), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT60), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n898), .A2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT119), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n944), .A3(new_n242), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n941), .B1(new_n841), .B2(new_n850), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT119), .B1(new_n946), .B2(new_n243), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n657), .B(KEYINPUT118), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n911), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n945), .A2(new_n947), .A3(new_n949), .A4(KEYINPUT61), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT61), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n898), .A2(new_n942), .A3(new_n948), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n912), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n946), .A2(new_n243), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n951), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n950), .A2(new_n955), .ZN(G66));
  INV_X1    g770(.A(new_n483), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n228), .B1(new_n957), .B2(new_n531), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT120), .Z(new_n959));
  OR2_X1    g773(.A1(new_n815), .A2(new_n822), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n961), .B2(G953), .ZN(new_n962));
  INV_X1    g776(.A(new_n902), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n963), .B1(G898), .B2(new_n228), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n962), .B(new_n964), .ZN(G69));
  AOI21_X1  g779(.A(new_n228), .B1(G227), .B2(G900), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n334), .B1(new_n314), .B2(new_n324), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n399), .B1(new_n401), .B2(new_n403), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n969), .A2(G953), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n675), .A2(new_n710), .A3(new_n739), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT62), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n706), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n706), .A2(new_n972), .ZN(new_n975));
  AOI21_X1  g789(.A(KEYINPUT121), .B1(new_n975), .B2(KEYINPUT62), .ZN(new_n976));
  INV_X1    g790(.A(KEYINPUT121), .ZN(new_n977));
  AOI211_X1 g791(.A(new_n977), .B(new_n973), .C1(new_n706), .C2(new_n972), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n800), .B(new_n974), .C1(new_n976), .C2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n789), .A2(new_n804), .ZN(new_n980));
  NOR3_X1   g794(.A1(new_n980), .A2(new_n679), .A3(new_n741), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n369), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n787), .A2(KEYINPUT122), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(KEYINPUT122), .B1(new_n787), .B2(new_n982), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n970), .B1(new_n979), .B2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n775), .A2(new_n609), .A3(new_n678), .ZN(new_n987));
  INV_X1    g801(.A(new_n691), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n885), .A2(new_n627), .A3(new_n988), .ZN(new_n989));
  OR3_X1    g803(.A1(new_n987), .A2(KEYINPUT125), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(KEYINPUT125), .B1(new_n987), .B2(new_n989), .ZN(new_n991));
  NAND4_X1  g805(.A1(new_n800), .A2(new_n990), .A3(new_n787), .A4(new_n991), .ZN(new_n992));
  OR3_X1    g806(.A1(new_n752), .A2(new_n971), .A3(new_n765), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n228), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n670), .A2(G953), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT124), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n994), .A2(new_n969), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n986), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n966), .B1(new_n998), .B2(KEYINPUT123), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT123), .ZN(new_n1000));
  INV_X1    g814(.A(new_n966), .ZN(new_n1001));
  AOI211_X1 g815(.A(new_n1000), .B(new_n1001), .C1(new_n986), .C2(new_n997), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n999), .A2(new_n1002), .ZN(G72));
  NAND2_X1  g817(.A1(G472), .A2(G902), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1004), .B(KEYINPUT63), .Z(new_n1005));
  NOR3_X1   g819(.A1(new_n357), .A2(KEYINPUT126), .A3(new_n252), .ZN(new_n1006));
  OAI21_X1  g820(.A(KEYINPUT126), .B1(new_n357), .B2(new_n252), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1007), .B1(new_n331), .B2(new_n332), .ZN(new_n1008));
  OAI221_X1 g822(.A(new_n1005), .B1(new_n1006), .B2(new_n1008), .C1(new_n831), .C2(new_n839), .ZN(new_n1009));
  NOR3_X1   g823(.A1(new_n992), .A2(new_n960), .A3(new_n993), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1005), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n363), .B(new_n357), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1009), .A2(new_n912), .A3(new_n1012), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n357), .A2(new_n363), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n979), .A2(new_n985), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1005), .B1(new_n1015), .B2(new_n960), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1013), .B1(new_n1014), .B2(new_n1016), .ZN(G57));
endmodule


