

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U556 ( .A(n749), .ZN(n727) );
  AND2_X1 U557 ( .A1(n843), .A2(n842), .ZN(n844) );
  OR2_X1 U558 ( .A1(n828), .A2(n827), .ZN(n843) );
  NOR2_X1 U559 ( .A1(n766), .A2(n765), .ZN(n823) );
  XNOR2_X1 U560 ( .A(n734), .B(n733), .ZN(n825) );
  BUF_X2 U561 ( .A(n580), .Z(n523) );
  INV_X1 U562 ( .A(n825), .ZN(n770) );
  XNOR2_X1 U563 ( .A(n748), .B(n747), .ZN(n755) );
  AND2_X1 U564 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U565 ( .A1(G543), .A2(G651), .ZN(n658) );
  NAND2_X1 U566 ( .A1(n826), .A2(n825), .ZN(n524) );
  AND2_X1 U567 ( .A1(n584), .A2(n583), .ZN(n525) );
  XNOR2_X1 U568 ( .A(n594), .B(KEYINPUT13), .ZN(n526) );
  OR2_X1 U569 ( .A1(n823), .A2(n822), .ZN(n527) );
  XNOR2_X1 U570 ( .A(KEYINPUT94), .B(KEYINPUT30), .ZN(n737) );
  INV_X1 U571 ( .A(KEYINPUT97), .ZN(n747) );
  INV_X1 U572 ( .A(G1966), .ZN(n735) );
  AND2_X1 U573 ( .A1(n825), .A2(n735), .ZN(n763) );
  NAND2_X1 U574 ( .A1(G160), .A2(G40), .ZN(n787) );
  INV_X1 U575 ( .A(n992), .ZN(n769) );
  INV_X1 U576 ( .A(KEYINPUT86), .ZN(n733) );
  NOR2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  NOR2_X1 U578 ( .A1(G651), .A2(n670), .ZN(n664) );
  XOR2_X1 U579 ( .A(G543), .B(KEYINPUT0), .Z(n670) );
  AND2_X1 U580 ( .A1(n525), .A2(n585), .ZN(n586) );
  NOR2_X2 U581 ( .A1(n537), .A2(n536), .ZN(G160) );
  INV_X1 U582 ( .A(G2104), .ZN(n528) );
  NOR2_X1 U583 ( .A1(n528), .A2(G2105), .ZN(n581) );
  NAND2_X1 U584 ( .A1(G101), .A2(n581), .ZN(n529) );
  XNOR2_X1 U585 ( .A(n529), .B(KEYINPUT23), .ZN(n530) );
  XNOR2_X1 U586 ( .A(n530), .B(KEYINPUT65), .ZN(n533) );
  XOR2_X1 U587 ( .A(KEYINPUT17), .B(n531), .Z(n580) );
  NAND2_X1 U588 ( .A1(G137), .A2(n523), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n533), .A2(n532), .ZN(n537) );
  AND2_X1 U590 ( .A1(n528), .A2(G2105), .ZN(n907) );
  NAND2_X1 U591 ( .A1(G125), .A2(n907), .ZN(n535) );
  AND2_X1 U592 ( .A1(G2104), .A2(G2105), .ZN(n908) );
  NAND2_X1 U593 ( .A1(G113), .A2(n908), .ZN(n534) );
  NAND2_X1 U594 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U595 ( .A1(n658), .A2(G89), .ZN(n538) );
  XNOR2_X1 U596 ( .A(n538), .B(KEYINPUT4), .ZN(n541) );
  INV_X1 U597 ( .A(G651), .ZN(n543) );
  OR2_X1 U598 ( .A1(n543), .A2(n670), .ZN(n539) );
  XOR2_X2 U599 ( .A(KEYINPUT66), .B(n539), .Z(n653) );
  NAND2_X1 U600 ( .A1(G76), .A2(n653), .ZN(n540) );
  NAND2_X1 U601 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U602 ( .A(n542), .B(KEYINPUT5), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G51), .A2(n664), .ZN(n546) );
  NOR2_X1 U604 ( .A1(G543), .A2(n543), .ZN(n544) );
  XOR2_X1 U605 ( .A(KEYINPUT1), .B(n544), .Z(n668) );
  NAND2_X1 U606 ( .A1(G63), .A2(n668), .ZN(n545) );
  NAND2_X1 U607 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U608 ( .A(KEYINPUT6), .B(n547), .Z(n548) );
  NAND2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U610 ( .A(n550), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U611 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U612 ( .A1(G85), .A2(n658), .ZN(n552) );
  NAND2_X1 U613 ( .A1(G72), .A2(n653), .ZN(n551) );
  NAND2_X1 U614 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U615 ( .A1(G47), .A2(n664), .ZN(n554) );
  NAND2_X1 U616 ( .A1(G60), .A2(n668), .ZN(n553) );
  NAND2_X1 U617 ( .A1(n554), .A2(n553), .ZN(n555) );
  OR2_X1 U618 ( .A1(n556), .A2(n555), .ZN(G290) );
  XOR2_X1 U619 ( .A(KEYINPUT106), .B(G2446), .Z(n558) );
  XNOR2_X1 U620 ( .A(G1341), .B(G1348), .ZN(n557) );
  XNOR2_X1 U621 ( .A(n558), .B(n557), .ZN(n570) );
  XOR2_X1 U622 ( .A(KEYINPUT105), .B(G2438), .Z(n560) );
  XNOR2_X1 U623 ( .A(KEYINPUT102), .B(KEYINPUT103), .ZN(n559) );
  XNOR2_X1 U624 ( .A(n560), .B(n559), .ZN(n568) );
  XOR2_X1 U625 ( .A(KEYINPUT107), .B(G2427), .Z(n562) );
  XNOR2_X1 U626 ( .A(G2454), .B(KEYINPUT104), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(n566) );
  XOR2_X1 U628 ( .A(G2451), .B(G2430), .Z(n564) );
  XNOR2_X1 U629 ( .A(G2443), .B(G2435), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(n566), .B(n565), .Z(n567) );
  XNOR2_X1 U632 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U633 ( .A(n570), .B(n569), .ZN(n571) );
  AND2_X1 U634 ( .A1(n571), .A2(G14), .ZN(G401) );
  NAND2_X1 U635 ( .A1(G52), .A2(n664), .ZN(n573) );
  NAND2_X1 U636 ( .A1(G64), .A2(n668), .ZN(n572) );
  NAND2_X1 U637 ( .A1(n573), .A2(n572), .ZN(n579) );
  NAND2_X1 U638 ( .A1(n658), .A2(G90), .ZN(n574) );
  XOR2_X1 U639 ( .A(KEYINPUT67), .B(n574), .Z(n576) );
  NAND2_X1 U640 ( .A1(G77), .A2(n653), .ZN(n575) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(KEYINPUT9), .B(n577), .Z(n578) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(G171) );
  AND2_X1 U644 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U645 ( .A(G57), .ZN(G237) );
  INV_X1 U646 ( .A(G132), .ZN(G219) );
  INV_X1 U647 ( .A(G82), .ZN(G220) );
  NAND2_X1 U648 ( .A1(n523), .A2(G138), .ZN(n587) );
  INV_X1 U649 ( .A(n581), .ZN(n582) );
  INV_X2 U650 ( .A(n582), .ZN(n912) );
  NAND2_X1 U651 ( .A1(G102), .A2(n912), .ZN(n584) );
  NAND2_X1 U652 ( .A1(G114), .A2(n908), .ZN(n583) );
  NAND2_X1 U653 ( .A1(G126), .A2(n907), .ZN(n585) );
  NAND2_X1 U654 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U655 ( .A(n588), .B(KEYINPUT79), .ZN(G164) );
  NAND2_X1 U656 ( .A1(G7), .A2(G661), .ZN(n589) );
  XNOR2_X1 U657 ( .A(n589), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U658 ( .A(G223), .ZN(n847) );
  NAND2_X1 U659 ( .A1(n847), .A2(G567), .ZN(n590) );
  XOR2_X1 U660 ( .A(KEYINPUT11), .B(n590), .Z(G234) );
  XOR2_X1 U661 ( .A(G860), .B(KEYINPUT71), .Z(n622) );
  NAND2_X1 U662 ( .A1(n658), .A2(G81), .ZN(n591) );
  XNOR2_X1 U663 ( .A(n591), .B(KEYINPUT12), .ZN(n593) );
  NAND2_X1 U664 ( .A1(G68), .A2(n653), .ZN(n592) );
  NAND2_X1 U665 ( .A1(n593), .A2(n592), .ZN(n594) );
  NAND2_X1 U666 ( .A1(G43), .A2(n664), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n526), .A2(n595), .ZN(n598) );
  NAND2_X1 U668 ( .A1(n668), .A2(G56), .ZN(n596) );
  XOR2_X1 U669 ( .A(KEYINPUT14), .B(n596), .Z(n597) );
  NOR2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n599) );
  XOR2_X2 U671 ( .A(KEYINPUT70), .B(n599), .Z(n998) );
  INV_X1 U672 ( .A(n998), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n622), .A2(n600), .ZN(G153) );
  INV_X1 U674 ( .A(G171), .ZN(G301) );
  INV_X1 U675 ( .A(G868), .ZN(n683) );
  NOR2_X1 U676 ( .A1(G301), .A2(n683), .ZN(n609) );
  NAND2_X1 U677 ( .A1(G92), .A2(n658), .ZN(n602) );
  NAND2_X1 U678 ( .A1(G79), .A2(n653), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U680 ( .A1(G54), .A2(n664), .ZN(n604) );
  NAND2_X1 U681 ( .A1(G66), .A2(n668), .ZN(n603) );
  NAND2_X1 U682 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U683 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U684 ( .A(KEYINPUT15), .B(n607), .Z(n991) );
  INV_X1 U685 ( .A(n991), .ZN(n624) );
  NOR2_X1 U686 ( .A1(G868), .A2(n624), .ZN(n608) );
  NOR2_X1 U687 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U688 ( .A(KEYINPUT72), .B(n610), .ZN(G284) );
  NAND2_X1 U689 ( .A1(G53), .A2(n664), .ZN(n612) );
  NAND2_X1 U690 ( .A1(G65), .A2(n668), .ZN(n611) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U692 ( .A(KEYINPUT69), .B(n613), .ZN(n618) );
  NAND2_X1 U693 ( .A1(G91), .A2(n658), .ZN(n615) );
  NAND2_X1 U694 ( .A1(G78), .A2(n653), .ZN(n614) );
  NAND2_X1 U695 ( .A1(n615), .A2(n614), .ZN(n616) );
  XOR2_X1 U696 ( .A(KEYINPUT68), .B(n616), .Z(n617) );
  NAND2_X1 U697 ( .A1(n618), .A2(n617), .ZN(G299) );
  NOR2_X1 U698 ( .A1(G286), .A2(n683), .ZN(n620) );
  NOR2_X1 U699 ( .A1(G868), .A2(G299), .ZN(n619) );
  NOR2_X1 U700 ( .A1(n620), .A2(n619), .ZN(G297) );
  INV_X1 U701 ( .A(G559), .ZN(n621) );
  NOR2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U704 ( .A(n625), .B(KEYINPUT73), .ZN(n626) );
  XNOR2_X1 U705 ( .A(n626), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U706 ( .A1(n998), .A2(G868), .ZN(n629) );
  NAND2_X1 U707 ( .A1(G868), .A2(n991), .ZN(n627) );
  NOR2_X1 U708 ( .A1(G559), .A2(n627), .ZN(n628) );
  NOR2_X1 U709 ( .A1(n629), .A2(n628), .ZN(G282) );
  NAND2_X1 U710 ( .A1(n907), .A2(G123), .ZN(n630) );
  XNOR2_X1 U711 ( .A(n630), .B(KEYINPUT18), .ZN(n632) );
  NAND2_X1 U712 ( .A1(G111), .A2(n908), .ZN(n631) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U714 ( .A1(G99), .A2(n912), .ZN(n634) );
  NAND2_X1 U715 ( .A1(G135), .A2(n523), .ZN(n633) );
  NAND2_X1 U716 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U717 ( .A1(n636), .A2(n635), .ZN(n944) );
  XNOR2_X1 U718 ( .A(G2096), .B(n944), .ZN(n638) );
  INV_X1 U719 ( .A(G2100), .ZN(n637) );
  NAND2_X1 U720 ( .A1(n638), .A2(n637), .ZN(G156) );
  NAND2_X1 U721 ( .A1(G559), .A2(n991), .ZN(n639) );
  XNOR2_X1 U722 ( .A(n639), .B(n998), .ZN(n680) );
  NOR2_X1 U723 ( .A1(G860), .A2(n680), .ZN(n646) );
  NAND2_X1 U724 ( .A1(G93), .A2(n658), .ZN(n641) );
  NAND2_X1 U725 ( .A1(G80), .A2(n653), .ZN(n640) );
  NAND2_X1 U726 ( .A1(n641), .A2(n640), .ZN(n645) );
  NAND2_X1 U727 ( .A1(G55), .A2(n664), .ZN(n643) );
  NAND2_X1 U728 ( .A1(G67), .A2(n668), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n643), .A2(n642), .ZN(n644) );
  OR2_X1 U730 ( .A1(n645), .A2(n644), .ZN(n682) );
  XOR2_X1 U731 ( .A(n646), .B(n682), .Z(G145) );
  NAND2_X1 U732 ( .A1(G88), .A2(n658), .ZN(n648) );
  NAND2_X1 U733 ( .A1(G75), .A2(n653), .ZN(n647) );
  NAND2_X1 U734 ( .A1(n648), .A2(n647), .ZN(n652) );
  NAND2_X1 U735 ( .A1(G50), .A2(n664), .ZN(n650) );
  NAND2_X1 U736 ( .A1(G62), .A2(n668), .ZN(n649) );
  NAND2_X1 U737 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U738 ( .A1(n652), .A2(n651), .ZN(G166) );
  NAND2_X1 U739 ( .A1(G73), .A2(n653), .ZN(n655) );
  XNOR2_X1 U740 ( .A(KEYINPUT2), .B(KEYINPUT76), .ZN(n654) );
  XNOR2_X1 U741 ( .A(n655), .B(n654), .ZN(n663) );
  NAND2_X1 U742 ( .A1(G48), .A2(n664), .ZN(n657) );
  NAND2_X1 U743 ( .A1(G61), .A2(n668), .ZN(n656) );
  NAND2_X1 U744 ( .A1(n657), .A2(n656), .ZN(n661) );
  NAND2_X1 U745 ( .A1(G86), .A2(n658), .ZN(n659) );
  XNOR2_X1 U746 ( .A(KEYINPUT75), .B(n659), .ZN(n660) );
  NOR2_X1 U747 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U748 ( .A1(n663), .A2(n662), .ZN(G305) );
  NAND2_X1 U749 ( .A1(G49), .A2(n664), .ZN(n666) );
  NAND2_X1 U750 ( .A1(G74), .A2(G651), .ZN(n665) );
  NAND2_X1 U751 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U752 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U753 ( .A(n669), .B(KEYINPUT74), .ZN(n672) );
  NAND2_X1 U754 ( .A1(G87), .A2(n670), .ZN(n671) );
  NAND2_X1 U755 ( .A1(n672), .A2(n671), .ZN(G288) );
  XOR2_X1 U756 ( .A(KEYINPUT77), .B(KEYINPUT19), .Z(n674) );
  XNOR2_X1 U757 ( .A(G166), .B(KEYINPUT78), .ZN(n673) );
  XNOR2_X1 U758 ( .A(n674), .B(n673), .ZN(n677) );
  INV_X1 U759 ( .A(G299), .ZN(n718) );
  XNOR2_X1 U760 ( .A(n718), .B(G305), .ZN(n675) );
  XNOR2_X1 U761 ( .A(n675), .B(G288), .ZN(n676) );
  XNOR2_X1 U762 ( .A(n677), .B(n676), .ZN(n679) );
  XOR2_X1 U763 ( .A(G290), .B(n682), .Z(n678) );
  XNOR2_X1 U764 ( .A(n679), .B(n678), .ZN(n856) );
  XNOR2_X1 U765 ( .A(n680), .B(n856), .ZN(n681) );
  NAND2_X1 U766 ( .A1(n681), .A2(G868), .ZN(n685) );
  NAND2_X1 U767 ( .A1(n683), .A2(n682), .ZN(n684) );
  NAND2_X1 U768 ( .A1(n685), .A2(n684), .ZN(G295) );
  NAND2_X1 U769 ( .A1(G2078), .A2(G2084), .ZN(n686) );
  XOR2_X1 U770 ( .A(KEYINPUT20), .B(n686), .Z(n687) );
  NAND2_X1 U771 ( .A1(G2090), .A2(n687), .ZN(n688) );
  XNOR2_X1 U772 ( .A(KEYINPUT21), .B(n688), .ZN(n689) );
  NAND2_X1 U773 ( .A1(n689), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U774 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U775 ( .A1(G220), .A2(G219), .ZN(n690) );
  XOR2_X1 U776 ( .A(KEYINPUT22), .B(n690), .Z(n691) );
  NOR2_X1 U777 ( .A1(G218), .A2(n691), .ZN(n692) );
  NAND2_X1 U778 ( .A1(G96), .A2(n692), .ZN(n854) );
  NAND2_X1 U779 ( .A1(n854), .A2(G2106), .ZN(n696) );
  NAND2_X1 U780 ( .A1(G69), .A2(G120), .ZN(n693) );
  NOR2_X1 U781 ( .A1(G237), .A2(n693), .ZN(n694) );
  NAND2_X1 U782 ( .A1(G108), .A2(n694), .ZN(n855) );
  NAND2_X1 U783 ( .A1(n855), .A2(G567), .ZN(n695) );
  NAND2_X1 U784 ( .A1(n696), .A2(n695), .ZN(n929) );
  NAND2_X1 U785 ( .A1(G483), .A2(G661), .ZN(n697) );
  NOR2_X1 U786 ( .A1(n929), .A2(n697), .ZN(n852) );
  NAND2_X1 U787 ( .A1(n852), .A2(G36), .ZN(G176) );
  INV_X1 U788 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U789 ( .A(G1981), .B(G305), .ZN(n983) );
  INV_X1 U790 ( .A(KEYINPUT32), .ZN(n758) );
  XNOR2_X1 U791 ( .A(KEYINPUT85), .B(n787), .ZN(n698) );
  NOR2_X1 U792 ( .A1(G164), .A2(G1384), .ZN(n788) );
  NAND2_X1 U793 ( .A1(n698), .A2(n788), .ZN(n749) );
  AND2_X1 U794 ( .A1(n727), .A2(G1996), .ZN(n700) );
  XOR2_X1 U795 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n699) );
  XNOR2_X1 U796 ( .A(n700), .B(n699), .ZN(n702) );
  NAND2_X1 U797 ( .A1(n749), .A2(G1341), .ZN(n701) );
  NAND2_X1 U798 ( .A1(n702), .A2(n701), .ZN(n703) );
  NOR2_X1 U799 ( .A1(n998), .A2(n703), .ZN(n704) );
  OR2_X1 U800 ( .A1(n991), .A2(n704), .ZN(n711) );
  NAND2_X1 U801 ( .A1(n991), .A2(n704), .ZN(n709) );
  AND2_X1 U802 ( .A1(n749), .A2(G1348), .ZN(n705) );
  XNOR2_X1 U803 ( .A(n705), .B(KEYINPUT93), .ZN(n707) );
  NAND2_X1 U804 ( .A1(n727), .A2(G2067), .ZN(n706) );
  NAND2_X1 U805 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U806 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U807 ( .A1(n711), .A2(n710), .ZN(n717) );
  XOR2_X1 U808 ( .A(KEYINPUT91), .B(KEYINPUT27), .Z(n713) );
  NAND2_X1 U809 ( .A1(G2072), .A2(n727), .ZN(n712) );
  XNOR2_X1 U810 ( .A(n713), .B(n712), .ZN(n715) );
  INV_X1 U811 ( .A(G1956), .ZN(n1005) );
  NOR2_X1 U812 ( .A1(n727), .A2(n1005), .ZN(n714) );
  NOR2_X1 U813 ( .A1(n715), .A2(n714), .ZN(n719) );
  NAND2_X1 U814 ( .A1(n719), .A2(n718), .ZN(n716) );
  NAND2_X1 U815 ( .A1(n717), .A2(n716), .ZN(n723) );
  NOR2_X1 U816 ( .A1(n719), .A2(n718), .ZN(n721) );
  XOR2_X1 U817 ( .A(KEYINPUT28), .B(KEYINPUT92), .Z(n720) );
  XNOR2_X1 U818 ( .A(n721), .B(n720), .ZN(n722) );
  NAND2_X1 U819 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U820 ( .A(KEYINPUT29), .B(n724), .ZN(n732) );
  XOR2_X1 U821 ( .A(G2078), .B(KEYINPUT25), .Z(n725) );
  XNOR2_X1 U822 ( .A(KEYINPUT88), .B(n725), .ZN(n961) );
  NOR2_X1 U823 ( .A1(n749), .A2(n961), .ZN(n726) );
  XOR2_X1 U824 ( .A(KEYINPUT89), .B(n726), .Z(n729) );
  NOR2_X1 U825 ( .A1(n727), .A2(G1961), .ZN(n728) );
  NOR2_X1 U826 ( .A1(n729), .A2(n728), .ZN(n740) );
  NOR2_X1 U827 ( .A1(n740), .A2(G301), .ZN(n730) );
  XNOR2_X1 U828 ( .A(n730), .B(KEYINPUT90), .ZN(n731) );
  NOR2_X1 U829 ( .A1(n732), .A2(n731), .ZN(n745) );
  NAND2_X1 U830 ( .A1(n749), .A2(G8), .ZN(n734) );
  NOR2_X1 U831 ( .A1(G2084), .A2(n749), .ZN(n760) );
  NOR2_X1 U832 ( .A1(n763), .A2(n760), .ZN(n736) );
  NAND2_X1 U833 ( .A1(n736), .A2(G8), .ZN(n738) );
  XNOR2_X1 U834 ( .A(n738), .B(n737), .ZN(n739) );
  NOR2_X1 U835 ( .A1(G168), .A2(n739), .ZN(n742) );
  AND2_X1 U836 ( .A1(G301), .A2(n740), .ZN(n741) );
  NOR2_X1 U837 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U838 ( .A(n743), .B(KEYINPUT31), .ZN(n744) );
  NOR2_X1 U839 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U840 ( .A(n746), .B(KEYINPUT95), .ZN(n759) );
  NAND2_X1 U841 ( .A1(n759), .A2(G286), .ZN(n748) );
  NOR2_X1 U842 ( .A1(G2090), .A2(n749), .ZN(n750) );
  XNOR2_X1 U843 ( .A(n750), .B(KEYINPUT98), .ZN(n752) );
  NOR2_X1 U844 ( .A1(n770), .A2(G1971), .ZN(n751) );
  NOR2_X1 U845 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U846 ( .A1(G303), .A2(n753), .ZN(n754) );
  NAND2_X1 U847 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U848 ( .A1(n756), .A2(G8), .ZN(n757) );
  XNOR2_X1 U849 ( .A(n758), .B(n757), .ZN(n766) );
  NAND2_X1 U850 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U851 ( .A1(n759), .A2(n761), .ZN(n762) );
  NOR2_X1 U852 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U853 ( .A(n764), .B(KEYINPUT96), .ZN(n765) );
  INV_X1 U854 ( .A(n823), .ZN(n768) );
  NOR2_X1 U855 ( .A1(G1976), .A2(G288), .ZN(n775) );
  NOR2_X1 U856 ( .A1(G1971), .A2(G303), .ZN(n767) );
  NOR2_X1 U857 ( .A1(n775), .A2(n767), .ZN(n986) );
  NAND2_X1 U858 ( .A1(n768), .A2(n986), .ZN(n772) );
  NAND2_X1 U859 ( .A1(G1976), .A2(G288), .ZN(n992) );
  NOR2_X1 U860 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U861 ( .A1(KEYINPUT33), .A2(n773), .ZN(n774) );
  NOR2_X1 U862 ( .A1(n983), .A2(n774), .ZN(n813) );
  AND2_X1 U863 ( .A1(n775), .A2(KEYINPUT33), .ZN(n776) );
  NAND2_X1 U864 ( .A1(n776), .A2(n825), .ZN(n811) );
  XOR2_X1 U865 ( .A(G1986), .B(G290), .Z(n985) );
  NAND2_X1 U866 ( .A1(n908), .A2(G116), .ZN(n777) );
  XOR2_X1 U867 ( .A(KEYINPUT81), .B(n777), .Z(n779) );
  NAND2_X1 U868 ( .A1(n907), .A2(G128), .ZN(n778) );
  NAND2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U870 ( .A(n780), .B(KEYINPUT35), .ZN(n785) );
  NAND2_X1 U871 ( .A1(G104), .A2(n912), .ZN(n782) );
  NAND2_X1 U872 ( .A1(G140), .A2(n523), .ZN(n781) );
  NAND2_X1 U873 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U874 ( .A(KEYINPUT34), .B(n783), .Z(n784) );
  NAND2_X1 U875 ( .A1(n785), .A2(n784), .ZN(n786) );
  XNOR2_X1 U876 ( .A(n786), .B(KEYINPUT36), .ZN(n920) );
  XOR2_X1 U877 ( .A(G2067), .B(KEYINPUT37), .Z(n829) );
  NAND2_X1 U878 ( .A1(n920), .A2(n829), .ZN(n936) );
  NAND2_X1 U879 ( .A1(n985), .A2(n936), .ZN(n790) );
  NOR2_X1 U880 ( .A1(n788), .A2(n787), .ZN(n789) );
  XOR2_X1 U881 ( .A(KEYINPUT80), .B(n789), .Z(n840) );
  INV_X1 U882 ( .A(n840), .ZN(n808) );
  AND2_X1 U883 ( .A1(n790), .A2(n808), .ZN(n810) );
  NAND2_X1 U884 ( .A1(n912), .A2(G105), .ZN(n791) );
  XNOR2_X1 U885 ( .A(n791), .B(KEYINPUT38), .ZN(n793) );
  NAND2_X1 U886 ( .A1(G141), .A2(n523), .ZN(n792) );
  NAND2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n797) );
  NAND2_X1 U888 ( .A1(G129), .A2(n907), .ZN(n795) );
  NAND2_X1 U889 ( .A1(G117), .A2(n908), .ZN(n794) );
  NAND2_X1 U890 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U891 ( .A1(n797), .A2(n796), .ZN(n798) );
  XNOR2_X1 U892 ( .A(KEYINPUT83), .B(n798), .ZN(n899) );
  NAND2_X1 U893 ( .A1(G1996), .A2(n899), .ZN(n807) );
  NAND2_X1 U894 ( .A1(G95), .A2(n912), .ZN(n800) );
  NAND2_X1 U895 ( .A1(G131), .A2(n523), .ZN(n799) );
  NAND2_X1 U896 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U897 ( .A1(n907), .A2(G119), .ZN(n801) );
  XOR2_X1 U898 ( .A(KEYINPUT82), .B(n801), .Z(n802) );
  NOR2_X1 U899 ( .A1(n803), .A2(n802), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n908), .A2(G107), .ZN(n804) );
  NAND2_X1 U901 ( .A1(n805), .A2(n804), .ZN(n904) );
  NAND2_X1 U902 ( .A1(G1991), .A2(n904), .ZN(n806) );
  NAND2_X1 U903 ( .A1(n807), .A2(n806), .ZN(n951) );
  NAND2_X1 U904 ( .A1(n951), .A2(n808), .ZN(n809) );
  XOR2_X1 U905 ( .A(KEYINPUT84), .B(n809), .Z(n832) );
  NOR2_X1 U906 ( .A1(n810), .A2(n832), .ZN(n814) );
  AND2_X1 U907 ( .A1(n811), .A2(n814), .ZN(n812) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n845) );
  INV_X1 U909 ( .A(n814), .ZN(n828) );
  INV_X1 U910 ( .A(G8), .ZN(n817) );
  NOR2_X1 U911 ( .A1(G2090), .A2(G303), .ZN(n815) );
  XNOR2_X1 U912 ( .A(n815), .B(KEYINPUT99), .ZN(n816) );
  NOR2_X1 U913 ( .A1(n817), .A2(n816), .ZN(n821) );
  NOR2_X1 U914 ( .A1(G1981), .A2(G305), .ZN(n818) );
  XOR2_X1 U915 ( .A(n818), .B(KEYINPUT87), .Z(n819) );
  XNOR2_X1 U916 ( .A(KEYINPUT24), .B(n819), .ZN(n820) );
  AND2_X1 U917 ( .A1(n825), .A2(n820), .ZN(n824) );
  OR2_X1 U918 ( .A1(n821), .A2(n824), .ZN(n822) );
  INV_X1 U919 ( .A(n824), .ZN(n826) );
  NAND2_X1 U920 ( .A1(n527), .A2(n524), .ZN(n827) );
  NOR2_X1 U921 ( .A1(n920), .A2(n829), .ZN(n947) );
  INV_X1 U922 ( .A(n936), .ZN(n837) );
  NOR2_X1 U923 ( .A1(G1996), .A2(n899), .ZN(n939) );
  NOR2_X1 U924 ( .A1(G1986), .A2(G290), .ZN(n830) );
  NOR2_X1 U925 ( .A1(G1991), .A2(n904), .ZN(n945) );
  NOR2_X1 U926 ( .A1(n830), .A2(n945), .ZN(n831) );
  NOR2_X1 U927 ( .A1(n832), .A2(n831), .ZN(n833) );
  NOR2_X1 U928 ( .A1(n939), .A2(n833), .ZN(n834) );
  XOR2_X1 U929 ( .A(n834), .B(KEYINPUT100), .Z(n835) );
  XNOR2_X1 U930 ( .A(KEYINPUT39), .B(n835), .ZN(n836) );
  NOR2_X1 U931 ( .A1(n837), .A2(n836), .ZN(n838) );
  NOR2_X1 U932 ( .A1(n947), .A2(n838), .ZN(n839) );
  NOR2_X1 U933 ( .A1(n840), .A2(n839), .ZN(n841) );
  XNOR2_X1 U934 ( .A(KEYINPUT101), .B(n841), .ZN(n842) );
  NAND2_X1 U935 ( .A1(n845), .A2(n844), .ZN(n846) );
  XNOR2_X1 U936 ( .A(n846), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U937 ( .A1(G2106), .A2(n847), .ZN(G217) );
  NAND2_X1 U938 ( .A1(G15), .A2(G2), .ZN(n848) );
  XOR2_X1 U939 ( .A(KEYINPUT108), .B(n848), .Z(n849) );
  NAND2_X1 U940 ( .A1(n849), .A2(G661), .ZN(n850) );
  XOR2_X1 U941 ( .A(KEYINPUT109), .B(n850), .Z(G259) );
  NAND2_X1 U942 ( .A1(G3), .A2(G1), .ZN(n851) );
  XNOR2_X1 U943 ( .A(KEYINPUT110), .B(n851), .ZN(n853) );
  NAND2_X1 U944 ( .A1(n853), .A2(n852), .ZN(G188) );
  INV_X1 U946 ( .A(G120), .ZN(G236) );
  INV_X1 U947 ( .A(G96), .ZN(G221) );
  INV_X1 U948 ( .A(G69), .ZN(G235) );
  NOR2_X1 U949 ( .A1(n855), .A2(n854), .ZN(G325) );
  INV_X1 U950 ( .A(G325), .ZN(G261) );
  XOR2_X1 U951 ( .A(n856), .B(G286), .Z(n858) );
  XNOR2_X1 U952 ( .A(n991), .B(G171), .ZN(n857) );
  XNOR2_X1 U953 ( .A(n858), .B(n857), .ZN(n859) );
  XNOR2_X1 U954 ( .A(n859), .B(n998), .ZN(n860) );
  NOR2_X1 U955 ( .A1(G37), .A2(n860), .ZN(G397) );
  XOR2_X1 U956 ( .A(KEYINPUT41), .B(G1986), .Z(n862) );
  XNOR2_X1 U957 ( .A(G1996), .B(G1991), .ZN(n861) );
  XNOR2_X1 U958 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U959 ( .A(n863), .B(KEYINPUT115), .Z(n865) );
  XNOR2_X1 U960 ( .A(G1981), .B(G1966), .ZN(n864) );
  XNOR2_X1 U961 ( .A(n865), .B(n864), .ZN(n869) );
  XOR2_X1 U962 ( .A(G1976), .B(G1971), .Z(n867) );
  XNOR2_X1 U963 ( .A(G1956), .B(G1961), .ZN(n866) );
  XNOR2_X1 U964 ( .A(n867), .B(n866), .ZN(n868) );
  XOR2_X1 U965 ( .A(n869), .B(n868), .Z(n871) );
  XNOR2_X1 U966 ( .A(KEYINPUT114), .B(G2474), .ZN(n870) );
  XNOR2_X1 U967 ( .A(n871), .B(n870), .ZN(G229) );
  XNOR2_X1 U968 ( .A(G2067), .B(G2078), .ZN(n872) );
  XNOR2_X1 U969 ( .A(n872), .B(KEYINPUT42), .ZN(n882) );
  XOR2_X1 U970 ( .A(G2678), .B(KEYINPUT43), .Z(n874) );
  XNOR2_X1 U971 ( .A(KEYINPUT112), .B(G2096), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n874), .B(n873), .ZN(n878) );
  XOR2_X1 U973 ( .A(G2100), .B(G2090), .Z(n876) );
  XNOR2_X1 U974 ( .A(G2072), .B(G2084), .ZN(n875) );
  XNOR2_X1 U975 ( .A(n876), .B(n875), .ZN(n877) );
  XOR2_X1 U976 ( .A(n878), .B(n877), .Z(n880) );
  XNOR2_X1 U977 ( .A(KEYINPUT113), .B(KEYINPUT111), .ZN(n879) );
  XNOR2_X1 U978 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(G227) );
  NAND2_X1 U980 ( .A1(n907), .A2(G124), .ZN(n883) );
  XNOR2_X1 U981 ( .A(n883), .B(KEYINPUT44), .ZN(n885) );
  NAND2_X1 U982 ( .A1(G112), .A2(n908), .ZN(n884) );
  NAND2_X1 U983 ( .A1(n885), .A2(n884), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G100), .A2(n912), .ZN(n887) );
  NAND2_X1 U985 ( .A1(G136), .A2(n523), .ZN(n886) );
  NAND2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n888) );
  NOR2_X1 U987 ( .A1(n889), .A2(n888), .ZN(G162) );
  XOR2_X1 U988 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n891) );
  XNOR2_X1 U989 ( .A(n944), .B(KEYINPUT117), .ZN(n890) );
  XNOR2_X1 U990 ( .A(n891), .B(n890), .ZN(n903) );
  NAND2_X1 U991 ( .A1(G103), .A2(n912), .ZN(n893) );
  NAND2_X1 U992 ( .A1(G139), .A2(n523), .ZN(n892) );
  NAND2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n898) );
  NAND2_X1 U994 ( .A1(G127), .A2(n907), .ZN(n895) );
  NAND2_X1 U995 ( .A1(G115), .A2(n908), .ZN(n894) );
  NAND2_X1 U996 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U997 ( .A(KEYINPUT47), .B(n896), .Z(n897) );
  NOR2_X1 U998 ( .A1(n898), .A2(n897), .ZN(n930) );
  XNOR2_X1 U999 ( .A(G160), .B(n930), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n899), .B(G164), .ZN(n900) );
  XNOR2_X1 U1001 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n903), .B(n902), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n904), .B(G162), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n919) );
  NAND2_X1 U1005 ( .A1(G130), .A2(n907), .ZN(n910) );
  NAND2_X1 U1006 ( .A1(G118), .A2(n908), .ZN(n909) );
  NAND2_X1 U1007 ( .A1(n910), .A2(n909), .ZN(n917) );
  NAND2_X1 U1008 ( .A1(n523), .A2(G142), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(n911), .B(KEYINPUT116), .ZN(n914) );
  NAND2_X1 U1010 ( .A1(G106), .A2(n912), .ZN(n913) );
  NAND2_X1 U1011 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1012 ( .A(n915), .B(KEYINPUT45), .Z(n916) );
  NOR2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1014 ( .A(n919), .B(n918), .Z(n921) );
  XNOR2_X1 U1015 ( .A(n921), .B(n920), .ZN(n922) );
  NOR2_X1 U1016 ( .A1(G37), .A2(n922), .ZN(G395) );
  NOR2_X1 U1017 ( .A1(G401), .A2(n929), .ZN(n926) );
  NOR2_X1 U1018 ( .A1(G229), .A2(G227), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(KEYINPUT49), .B(n923), .ZN(n924) );
  NOR2_X1 U1020 ( .A1(G397), .A2(n924), .ZN(n925) );
  NAND2_X1 U1021 ( .A1(n926), .A2(n925), .ZN(n927) );
  NOR2_X1 U1022 ( .A1(n927), .A2(G395), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(n928), .B(KEYINPUT118), .ZN(G308) );
  INV_X1 U1024 ( .A(G308), .ZN(G225) );
  INV_X1 U1025 ( .A(n929), .ZN(G319) );
  INV_X1 U1026 ( .A(G108), .ZN(G238) );
  INV_X1 U1027 ( .A(KEYINPUT55), .ZN(n957) );
  XNOR2_X1 U1028 ( .A(G164), .B(G2078), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(G2072), .B(n930), .ZN(n931) );
  XNOR2_X1 U1030 ( .A(n931), .B(KEYINPUT120), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1032 ( .A(n934), .B(KEYINPUT50), .ZN(n935) );
  XNOR2_X1 U1033 ( .A(n935), .B(KEYINPUT121), .ZN(n937) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n943) );
  XNOR2_X1 U1035 ( .A(G2090), .B(G162), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(n938), .B(KEYINPUT119), .ZN(n940) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(KEYINPUT51), .B(n941), .ZN(n942) );
  NOR2_X1 U1039 ( .A1(n943), .A2(n942), .ZN(n953) );
  NOR2_X1 U1040 ( .A1(n945), .A2(n944), .ZN(n949) );
  XOR2_X1 U1041 ( .A(G2084), .B(G160), .Z(n946) );
  NOR2_X1 U1042 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n949), .A2(n948), .ZN(n950) );
  NOR2_X1 U1044 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1045 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1046 ( .A(KEYINPUT52), .B(n954), .ZN(n955) );
  XOR2_X1 U1047 ( .A(KEYINPUT122), .B(n955), .Z(n956) );
  NAND2_X1 U1048 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1049 ( .A1(n958), .A2(G29), .ZN(n1034) );
  XOR2_X1 U1050 ( .A(G29), .B(KEYINPUT126), .Z(n980) );
  XNOR2_X1 U1051 ( .A(G2072), .B(G33), .ZN(n960) );
  XNOR2_X1 U1052 ( .A(G2067), .B(G26), .ZN(n959) );
  NOR2_X1 U1053 ( .A1(n960), .A2(n959), .ZN(n965) );
  XNOR2_X1 U1054 ( .A(n961), .B(G27), .ZN(n963) );
  XNOR2_X1 U1055 ( .A(G32), .B(G1996), .ZN(n962) );
  NOR2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n964) );
  NAND2_X1 U1057 ( .A1(n965), .A2(n964), .ZN(n969) );
  XOR2_X1 U1058 ( .A(G1991), .B(G25), .Z(n966) );
  NAND2_X1 U1059 ( .A1(n966), .A2(G28), .ZN(n967) );
  XNOR2_X1 U1060 ( .A(KEYINPUT124), .B(n967), .ZN(n968) );
  NOR2_X1 U1061 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1062 ( .A(n970), .B(KEYINPUT53), .ZN(n971) );
  XNOR2_X1 U1063 ( .A(n971), .B(KEYINPUT125), .ZN(n974) );
  XOR2_X1 U1064 ( .A(G2084), .B(G34), .Z(n972) );
  XNOR2_X1 U1065 ( .A(KEYINPUT54), .B(n972), .ZN(n973) );
  NAND2_X1 U1066 ( .A1(n974), .A2(n973), .ZN(n977) );
  XOR2_X1 U1067 ( .A(KEYINPUT123), .B(G2090), .Z(n975) );
  XNOR2_X1 U1068 ( .A(G35), .B(n975), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(n978), .B(KEYINPUT55), .ZN(n979) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1072 ( .A1(G11), .A2(n981), .ZN(n1032) );
  XNOR2_X1 U1073 ( .A(G16), .B(KEYINPUT56), .ZN(n1004) );
  XOR2_X1 U1074 ( .A(G168), .B(G1966), .Z(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  XOR2_X1 U1076 ( .A(KEYINPUT57), .B(n984), .Z(n1002) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n988) );
  XNOR2_X1 U1078 ( .A(G1956), .B(G299), .ZN(n987) );
  NOR2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n997) );
  XNOR2_X1 U1080 ( .A(G171), .B(G1961), .ZN(n990) );
  NAND2_X1 U1081 ( .A1(G1971), .A2(G303), .ZN(n989) );
  NAND2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(n991), .B(G1348), .ZN(n993) );
  NAND2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n1000) );
  XNOR2_X1 U1087 ( .A(G1341), .B(n998), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1089 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1090 ( .A1(n1004), .A2(n1003), .ZN(n1030) );
  INV_X1 U1091 ( .A(G16), .ZN(n1028) );
  XNOR2_X1 U1092 ( .A(G20), .B(n1005), .ZN(n1009) );
  XNOR2_X1 U1093 ( .A(G1981), .B(G6), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(G1341), .B(G19), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NAND2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1012) );
  XOR2_X1 U1097 ( .A(KEYINPUT59), .B(G1348), .Z(n1010) );
  XNOR2_X1 U1098 ( .A(G4), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(KEYINPUT60), .B(n1013), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(G1966), .B(G21), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(G1961), .B(G5), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1104 ( .A1(n1017), .A2(n1016), .ZN(n1025) );
  XNOR2_X1 U1105 ( .A(G1976), .B(G23), .ZN(n1019) );
  XNOR2_X1 U1106 ( .A(G1986), .B(G24), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(G1971), .B(KEYINPUT127), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(n1020), .B(G22), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1111 ( .A(KEYINPUT58), .B(n1023), .ZN(n1024) );
  NOR2_X1 U1112 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1113 ( .A(KEYINPUT61), .B(n1026), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1035), .Z(G311) );
  INV_X1 U1119 ( .A(G311), .ZN(G150) );
endmodule

