//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 1 1 1 0 1 1 0 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n536,
    new_n537, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n550, new_n551, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n594, new_n595,
    new_n598, new_n600, new_n601, new_n602, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1178,
    new_n1179, new_n1180;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  AND2_X1   g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G101), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G137), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT65), .B(G2105), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT65), .A2(G2105), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n468), .A2(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(new_n471), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n479), .A2(G2105), .ZN(new_n481));
  AOI22_X1  g056(.A1(G124), .A2(new_n480), .B1(new_n481), .B2(G136), .ZN(new_n482));
  OAI221_X1 g057(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n471), .C2(G112), .ZN(new_n483));
  AND2_X1   g058(.A1(new_n482), .A2(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n485));
  INV_X1    g060(.A(G114), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g064(.A(G138), .B1(new_n464), .B2(new_n465), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT4), .B1(new_n490), .B2(new_n467), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n478), .A2(new_n471), .A3(new_n492), .A4(G138), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(G164));
  INV_X1    g069(.A(G651), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G62), .ZN(new_n501));
  OR2_X1    g076(.A1(new_n501), .A2(KEYINPUT66), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n501), .A2(KEYINPUT66), .B1(G75), .B2(G543), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n495), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n505), .A2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n506), .A2(new_n507), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n504), .A2(new_n510), .ZN(G166));
  NAND3_X1  g086(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n512), .B(KEYINPUT7), .ZN(new_n513));
  INV_X1    g088(.A(new_n506), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G89), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n500), .A2(G63), .A3(G651), .ZN(new_n516));
  INV_X1    g091(.A(G51), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n508), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g093(.A(new_n513), .B(new_n515), .C1(new_n518), .C2(KEYINPUT67), .ZN(new_n519));
  AND2_X1   g094(.A1(new_n518), .A2(KEYINPUT67), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(G168));
  AOI22_X1  g096(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n522), .A2(new_n495), .ZN(new_n523));
  INV_X1    g098(.A(G90), .ZN(new_n524));
  INV_X1    g099(.A(G52), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n506), .A2(new_n524), .B1(new_n508), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G171));
  AOI22_X1  g102(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n495), .ZN(new_n529));
  INV_X1    g104(.A(G81), .ZN(new_n530));
  INV_X1    g105(.A(G43), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n506), .A2(new_n530), .B1(new_n508), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n529), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G860), .ZN(G153));
  NAND4_X1  g109(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g110(.A1(G1), .A2(G3), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT8), .ZN(new_n537));
  NAND4_X1  g112(.A1(G319), .A2(G483), .A3(G661), .A4(new_n537), .ZN(G188));
  INV_X1    g113(.A(KEYINPUT68), .ZN(new_n539));
  NAND4_X1  g114(.A1(new_n505), .A2(new_n539), .A3(G53), .A4(G543), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT9), .ZN(new_n541));
  NAND2_X1  g116(.A1(G78), .A2(G543), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n498), .A2(new_n499), .ZN(new_n543));
  INV_X1    g118(.A(G65), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n545), .A2(G651), .B1(new_n514), .B2(G91), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT69), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n547), .B(new_n548), .ZN(G299));
  INV_X1    g124(.A(KEYINPUT70), .ZN(new_n550));
  XNOR2_X1  g125(.A(G171), .B(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(G301));
  INV_X1    g127(.A(G168), .ZN(G286));
  INV_X1    g128(.A(G166), .ZN(G303));
  NAND2_X1  g129(.A1(G74), .A2(G651), .ZN(new_n555));
  OAI211_X1 g130(.A(KEYINPUT71), .B(new_n555), .C1(new_n543), .C2(new_n495), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT71), .ZN(new_n557));
  OAI211_X1 g132(.A(new_n557), .B(G651), .C1(new_n500), .C2(G74), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n505), .A2(G49), .A3(G543), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n500), .A2(new_n505), .A3(G87), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n556), .A2(new_n558), .A3(new_n559), .A4(new_n560), .ZN(G288));
  NAND2_X1  g136(.A1(new_n514), .A2(G86), .ZN(new_n562));
  AND2_X1   g137(.A1(new_n505), .A2(G543), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G48), .ZN(new_n564));
  NAND2_X1  g139(.A1(G73), .A2(G543), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT72), .ZN(new_n566));
  INV_X1    g141(.A(G61), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n567), .B1(new_n498), .B2(new_n499), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n562), .A2(new_n564), .A3(new_n569), .ZN(G305));
  AOI22_X1  g145(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n571), .A2(new_n495), .ZN(new_n572));
  INV_X1    g147(.A(G85), .ZN(new_n573));
  INV_X1    g148(.A(G47), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n506), .A2(new_n573), .B1(new_n508), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G290));
  NAND2_X1  g152(.A1(G79), .A2(G543), .ZN(new_n578));
  INV_X1    g153(.A(G66), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n543), .B2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n580), .A2(G651), .B1(new_n563), .B2(G54), .ZN(new_n581));
  XOR2_X1   g156(.A(KEYINPUT74), .B(KEYINPUT10), .Z(new_n582));
  NAND3_X1  g157(.A1(new_n514), .A2(G92), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n582), .ZN(new_n584));
  INV_X1    g159(.A(G92), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n506), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n581), .A2(new_n583), .A3(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT73), .B1(new_n588), .B2(G868), .ZN(new_n589));
  INV_X1    g164(.A(G868), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n551), .A2(new_n590), .ZN(new_n591));
  MUX2_X1   g166(.A(new_n589), .B(KEYINPUT73), .S(new_n591), .Z(G284));
  MUX2_X1   g167(.A(new_n589), .B(KEYINPUT73), .S(new_n591), .Z(G321));
  NAND2_X1  g168(.A1(G286), .A2(G868), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n547), .B(KEYINPUT69), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(G868), .ZN(G297));
  OAI21_X1  g171(.A(new_n594), .B1(new_n595), .B2(G868), .ZN(G280));
  INV_X1    g172(.A(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n588), .B1(new_n598), .B2(G860), .ZN(G148));
  INV_X1    g174(.A(new_n533), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n600), .A2(new_n590), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n587), .A2(G559), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(new_n590), .ZN(G323));
  XNOR2_X1  g178(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g179(.A1(new_n478), .A2(new_n462), .ZN(new_n605));
  XOR2_X1   g180(.A(KEYINPUT75), .B(KEYINPUT12), .Z(new_n606));
  XNOR2_X1  g181(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2100), .ZN(new_n609));
  AOI22_X1  g184(.A1(G123), .A2(new_n480), .B1(new_n481), .B2(G135), .ZN(new_n610));
  OAI221_X1 g185(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n471), .C2(G111), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g187(.A(KEYINPUT76), .B(G2096), .Z(new_n613));
  XNOR2_X1  g188(.A(new_n612), .B(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n609), .A2(new_n614), .ZN(G156));
  XNOR2_X1  g190(.A(G2427), .B(G2438), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(G2430), .ZN(new_n617));
  XNOR2_X1  g192(.A(KEYINPUT15), .B(G2435), .ZN(new_n618));
  OR2_X1    g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n619), .A2(KEYINPUT14), .A3(new_n620), .ZN(new_n621));
  XNOR2_X1  g196(.A(G2443), .B(G2446), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G1341), .B(G1348), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(G2451), .B(G2454), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT16), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT77), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n625), .A2(new_n628), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(G14), .A3(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(new_n631), .ZN(G401));
  XOR2_X1   g207(.A(G2072), .B(G2078), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT17), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2067), .B(G2678), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  NOR2_X1   g211(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g212(.A(KEYINPUT78), .ZN(new_n638));
  XOR2_X1   g213(.A(G2084), .B(G2090), .Z(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(new_n636), .B2(new_n633), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n637), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(new_n638), .B2(new_n640), .ZN(new_n642));
  INV_X1    g217(.A(new_n633), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n643), .A2(new_n639), .A3(new_n635), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT18), .Z(new_n645));
  NAND3_X1  g220(.A1(new_n634), .A2(new_n639), .A3(new_n636), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n642), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2096), .B(G2100), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(G227));
  XOR2_X1   g224(.A(G1971), .B(G1976), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT19), .ZN(new_n651));
  XNOR2_X1  g226(.A(G1956), .B(G2474), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G1961), .B(G1966), .Z(new_n654));
  AND2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT20), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n653), .A2(new_n654), .ZN(new_n658));
  NOR3_X1   g233(.A1(new_n651), .A2(new_n655), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n659), .B1(new_n651), .B2(new_n658), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1991), .B(G1996), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n663), .B(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G1981), .B(G1986), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G229));
  INV_X1    g242(.A(G29), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(G32), .ZN(new_n669));
  NAND3_X1  g244(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT26), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n481), .A2(G141), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n462), .A2(G105), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI211_X1 g249(.A(new_n671), .B(new_n674), .C1(G129), .C2(new_n480), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n669), .B1(new_n675), .B2(new_n668), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT27), .B(G1996), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT83), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT24), .B(G34), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n680), .A2(new_n668), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT82), .Z(new_n682));
  INV_X1    g257(.A(G160), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n682), .B1(new_n683), .B2(new_n668), .ZN(new_n684));
  INV_X1    g259(.A(G2084), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G16), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n687), .A2(G19), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n533), .B2(new_n687), .ZN(new_n689));
  XOR2_X1   g264(.A(new_n689), .B(G1341), .Z(new_n690));
  NOR2_X1   g265(.A1(G171), .A2(new_n687), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G5), .B2(new_n687), .ZN(new_n692));
  INV_X1    g267(.A(G1961), .ZN(new_n693));
  AOI22_X1  g268(.A1(new_n692), .A2(new_n693), .B1(new_n685), .B2(new_n684), .ZN(new_n694));
  NAND4_X1  g269(.A1(new_n679), .A2(new_n686), .A3(new_n690), .A4(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(G29), .A2(G35), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n696), .B1(G162), .B2(G29), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(G2090), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT89), .B(KEYINPUT29), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n668), .A2(G26), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(KEYINPUT28), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n481), .A2(G140), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n480), .A2(G128), .ZN(new_n704));
  OAI221_X1 g279(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n471), .C2(G116), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n702), .B1(new_n706), .B2(G29), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(G2067), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n668), .A2(G27), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G164), .B2(new_n668), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(G2078), .Z(new_n711));
  NAND2_X1  g286(.A1(new_n588), .A2(G16), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G4), .B2(G16), .ZN(new_n713));
  INV_X1    g288(.A(G1348), .ZN(new_n714));
  OAI211_X1 g289(.A(new_n708), .B(new_n711), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n668), .A2(G33), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n471), .A2(G103), .A3(G2104), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n717), .B(KEYINPUT25), .Z(new_n718));
  NAND2_X1  g293(.A1(G115), .A2(G2104), .ZN(new_n719));
  INV_X1    g294(.A(G127), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(new_n479), .B2(new_n720), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n721), .A2(new_n467), .B1(new_n481), .B2(G139), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n718), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n716), .B1(new_n724), .B2(new_n668), .ZN(new_n725));
  AOI22_X1  g300(.A1(new_n713), .A2(new_n714), .B1(new_n725), .B2(G2072), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G2072), .B2(new_n725), .ZN(new_n727));
  NOR4_X1   g302(.A1(new_n695), .A2(new_n700), .A3(new_n715), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n687), .A2(G20), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT23), .Z(new_n730));
  AOI21_X1  g305(.A(new_n730), .B1(G299), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G1956), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n692), .A2(new_n693), .ZN(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT87), .Z(new_n735));
  NAND2_X1  g310(.A1(G168), .A2(G16), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT84), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n736), .B(new_n737), .C1(G16), .C2(G21), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n737), .B2(new_n736), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(G1966), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(G1966), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n612), .A2(new_n668), .ZN(new_n742));
  OR2_X1    g317(.A1(new_n742), .A2(KEYINPUT85), .ZN(new_n743));
  XOR2_X1   g318(.A(KEYINPUT31), .B(G11), .Z(new_n744));
  XOR2_X1   g319(.A(KEYINPUT86), .B(G28), .Z(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(KEYINPUT30), .ZN(new_n746));
  AOI21_X1  g321(.A(G29), .B1(new_n745), .B2(KEYINPUT30), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n744), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n743), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(KEYINPUT85), .B2(new_n742), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n735), .A2(new_n740), .A3(new_n741), .A4(new_n750), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n728), .B(new_n732), .C1(new_n733), .C2(new_n751), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n751), .A2(new_n733), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT36), .ZN(new_n756));
  OR2_X1    g331(.A1(G6), .A2(G16), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(G305), .B2(new_n687), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT32), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(G1981), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n687), .A2(G22), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(G166), .B2(new_n687), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G1971), .Z(new_n763));
  MUX2_X1   g338(.A(G23), .B(G288), .S(G16), .Z(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT33), .B(G1976), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n760), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT80), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  NAND3_X1  g345(.A1(new_n769), .A2(KEYINPUT34), .A3(new_n770), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT81), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(KEYINPUT34), .B1(new_n769), .B2(new_n770), .ZN(new_n774));
  OR2_X1    g349(.A1(G25), .A2(G29), .ZN(new_n775));
  OAI221_X1 g350(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n471), .C2(G107), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT79), .ZN(new_n777));
  AOI22_X1  g352(.A1(G119), .A2(new_n480), .B1(new_n481), .B2(G131), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n775), .B1(new_n779), .B2(new_n668), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT35), .B(G1991), .Z(new_n781));
  NOR2_X1   g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n687), .A2(G24), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n576), .B2(new_n687), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1986), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n774), .A2(new_n782), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n756), .B1(new_n773), .B2(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n773), .A2(new_n787), .A3(new_n756), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n755), .B1(new_n789), .B2(new_n790), .ZN(G311));
  INV_X1    g366(.A(new_n790), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n754), .B1(new_n792), .B2(new_n788), .ZN(G150));
  AOI22_X1  g368(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n794), .A2(new_n495), .ZN(new_n795));
  INV_X1    g370(.A(G93), .ZN(new_n796));
  INV_X1    g371(.A(G55), .ZN(new_n797));
  OAI22_X1  g372(.A1(new_n506), .A2(new_n796), .B1(new_n508), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(G860), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(KEYINPUT37), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n795), .A2(new_n798), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT91), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n799), .A2(KEYINPUT91), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n805), .A2(new_n533), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n600), .A2(new_n803), .A3(new_n804), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n588), .A2(G559), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT90), .B(KEYINPUT38), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n800), .B1(new_n814), .B2(KEYINPUT39), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n802), .B1(new_n815), .B2(new_n816), .ZN(G145));
  INV_X1    g392(.A(KEYINPUT40), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n779), .B(new_n607), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n481), .A2(G142), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT95), .Z(new_n821));
  NAND2_X1  g396(.A1(new_n480), .A2(G130), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n471), .A2(G118), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n821), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n819), .B(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT96), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n491), .A2(new_n493), .ZN(new_n829));
  NAND2_X1  g404(.A1(G126), .A2(G2105), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n830), .B1(new_n476), .B2(new_n477), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n461), .A2(G114), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(KEYINPUT93), .B1(new_n831), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n485), .A2(new_n488), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n829), .A2(new_n835), .A3(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n706), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n675), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n724), .A2(KEYINPUT94), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n724), .A2(KEYINPUT94), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n840), .B1(new_n841), .B2(new_n843), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n828), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n826), .A2(new_n827), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(G162), .B(G160), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(KEYINPUT92), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n849), .B(new_n612), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(G37), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n847), .A2(new_n850), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n818), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n854), .ZN(new_n856));
  NAND4_X1  g431(.A1(new_n856), .A2(KEYINPUT40), .A3(new_n852), .A4(new_n851), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n855), .A2(new_n857), .ZN(G395));
  INV_X1    g433(.A(KEYINPUT99), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT97), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n807), .A2(new_n808), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n602), .ZN(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(G299), .A2(new_n588), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n595), .A2(new_n587), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n860), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT41), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n864), .A2(new_n865), .A3(KEYINPUT41), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n862), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n867), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n860), .A3(new_n862), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n859), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n873), .A2(new_n859), .A3(new_n874), .ZN(new_n876));
  XNOR2_X1  g451(.A(G166), .B(G290), .ZN(new_n877));
  XOR2_X1   g452(.A(G305), .B(G288), .Z(new_n878));
  XOR2_X1   g453(.A(new_n877), .B(new_n878), .Z(new_n879));
  NOR3_X1   g454(.A1(new_n879), .A2(KEYINPUT98), .A3(KEYINPUT42), .ZN(new_n880));
  XOR2_X1   g455(.A(KEYINPUT98), .B(KEYINPUT42), .Z(new_n881));
  AOI21_X1  g456(.A(new_n880), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  AND3_X1   g457(.A1(new_n875), .A2(new_n876), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n875), .B1(new_n876), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g459(.A(G868), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n885), .B1(G868), .B2(new_n799), .ZN(G295));
  OAI21_X1  g461(.A(new_n885), .B1(G868), .B2(new_n799), .ZN(G331));
  NAND2_X1  g462(.A1(new_n551), .A2(G168), .ZN(new_n888));
  OR2_X1    g463(.A1(G168), .A2(G171), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(new_n809), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n861), .A2(new_n888), .A3(new_n889), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n871), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n891), .A2(new_n892), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(new_n866), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(KEYINPUT100), .A3(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n896), .A2(KEYINPUT100), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(KEYINPUT101), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT101), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n901), .A3(new_n898), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n900), .A2(new_n879), .A3(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(new_n879), .ZN(new_n904));
  AOI21_X1  g479(.A(G37), .B1(new_n899), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT43), .B1(new_n903), .B2(new_n905), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n895), .A2(new_n866), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT41), .B1(new_n864), .B2(new_n865), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n895), .B1(KEYINPUT102), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT102), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n869), .A2(new_n910), .A3(new_n870), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n907), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT103), .B1(new_n912), .B2(new_n904), .ZN(new_n913));
  INV_X1    g488(.A(new_n911), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n891), .B(new_n892), .C1(new_n869), .C2(new_n910), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n896), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n917), .A3(new_n879), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n913), .A2(new_n918), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n919), .A2(new_n905), .A3(KEYINPUT43), .ZN(new_n920));
  OAI21_X1  g495(.A(KEYINPUT44), .B1(new_n906), .B2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT43), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n903), .B2(new_n905), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n919), .A2(new_n905), .A3(new_n923), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n921), .A2(new_n926), .ZN(G397));
  XOR2_X1   g502(.A(KEYINPUT104), .B(G1384), .Z(new_n928));
  NAND2_X1  g503(.A1(new_n838), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT45), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(G160), .A2(G40), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G1996), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n935), .A3(new_n675), .ZN(new_n936));
  XOR2_X1   g511(.A(new_n936), .B(KEYINPUT105), .Z(new_n937));
  XOR2_X1   g512(.A(new_n706), .B(G2067), .Z(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT106), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n934), .B1(new_n939), .B2(new_n675), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n935), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n942), .A2(new_n777), .A3(new_n778), .A4(new_n781), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n706), .A2(G2067), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n934), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n779), .B(new_n781), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n942), .B1(new_n934), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(G1986), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n933), .A2(new_n948), .A3(new_n576), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n949), .B(KEYINPUT48), .Z(new_n950));
  NOR2_X1   g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n933), .A2(new_n935), .ZN(new_n952));
  XOR2_X1   g527(.A(new_n952), .B(KEYINPUT46), .Z(new_n953));
  NOR2_X1   g528(.A1(new_n940), .A2(new_n953), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n954), .B(KEYINPUT47), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n945), .A2(new_n951), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT114), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT9), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n540), .B(new_n958), .ZN(new_n959));
  AOI22_X1  g534(.A1(new_n500), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n960));
  INV_X1    g535(.A(G91), .ZN(new_n961));
  OAI22_X1  g536(.A1(new_n960), .A2(new_n495), .B1(new_n961), .B2(new_n506), .ZN(new_n962));
  OAI211_X1 g537(.A(new_n957), .B(KEYINPUT57), .C1(new_n959), .C2(new_n962), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n957), .A2(KEYINPUT57), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n957), .A2(KEYINPUT57), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n541), .A2(new_n546), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(new_n966), .ZN(new_n967));
  NOR2_X1   g542(.A1(G164), .A2(G1384), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT50), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n932), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n838), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT50), .ZN(new_n973));
  AOI21_X1  g548(.A(G1956), .B1(new_n970), .B2(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n491), .A2(new_n493), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n835), .A2(new_n837), .ZN(new_n976));
  OAI211_X1 g551(.A(KEYINPUT45), .B(new_n928), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n930), .B1(G164), .B2(G1384), .ZN(new_n978));
  INV_X1    g553(.A(G40), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n468), .A2(new_n474), .A3(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT56), .B(G2072), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n977), .A2(new_n978), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n967), .B1(new_n974), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n838), .A2(new_n971), .A3(new_n980), .ZN(new_n985));
  NOR2_X1   g560(.A1(new_n985), .A2(G2067), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT50), .B1(new_n838), .B2(new_n971), .ZN(new_n987));
  NOR3_X1   g562(.A1(G164), .A2(new_n969), .A3(G1384), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n980), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n986), .B1(new_n989), .B2(new_n714), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n984), .B1(new_n587), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1956), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n831), .A2(new_n834), .ZN(new_n993));
  INV_X1    g568(.A(G138), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n476), .B2(new_n477), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n492), .B1(new_n995), .B2(new_n471), .ZN(new_n996));
  NOR3_X1   g571(.A1(new_n490), .A2(new_n467), .A3(KEYINPUT4), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n993), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n998), .A2(new_n969), .A3(new_n971), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n980), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n969), .B1(new_n838), .B2(new_n971), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n992), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AND2_X1   g577(.A1(new_n963), .A2(new_n966), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n1003), .A3(new_n982), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n991), .A2(KEYINPUT115), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  AOI21_X1  g581(.A(KEYINPUT115), .B1(new_n991), .B2(new_n1004), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT61), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n974), .A2(new_n983), .A3(new_n967), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1003), .B1(new_n1002), .B2(new_n982), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT118), .ZN(new_n1013));
  NAND4_X1  g588(.A1(new_n977), .A2(new_n978), .A3(new_n935), .A4(new_n980), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT58), .B(G1341), .Z(new_n1015));
  NAND2_X1  g590(.A1(new_n985), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT117), .B1(new_n1017), .B2(new_n533), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT117), .ZN(new_n1019));
  AOI211_X1 g594(.A(new_n1019), .B(new_n600), .C1(new_n1014), .C2(new_n1016), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT59), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1022), .A2(KEYINPUT116), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1012), .A2(new_n1013), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  OAI22_X1  g599(.A1(new_n1018), .A2(new_n1020), .B1(KEYINPUT116), .B2(new_n1022), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n984), .A2(new_n1004), .A3(KEYINPUT61), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  OAI211_X1 g602(.A(KEYINPUT118), .B(new_n1009), .C1(new_n1010), .C2(new_n1011), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n1024), .A2(new_n1027), .A3(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n990), .A2(KEYINPUT60), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT60), .ZN(new_n1031));
  AOI211_X1 g606(.A(new_n1031), .B(new_n986), .C1(new_n989), .C2(new_n714), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n588), .B1(new_n1032), .B2(KEYINPUT119), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n990), .A2(KEYINPUT60), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT119), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1034), .A2(new_n1035), .A3(new_n587), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1032), .A2(KEYINPUT119), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1030), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1008), .B1(new_n1029), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(G286), .A2(G8), .ZN(new_n1041));
  INV_X1    g616(.A(G1966), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n998), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n980), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT45), .B1(new_n838), .B2(new_n971), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT112), .B(G2084), .Z(new_n1047));
  NOR2_X1   g622(.A1(new_n932), .A2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g623(.A(KEYINPUT113), .B(new_n1048), .C1(new_n987), .C2(new_n988), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n998), .A2(KEYINPUT50), .A3(new_n971), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n835), .A2(new_n837), .ZN(new_n1052));
  AOI21_X1  g627(.A(G1384), .B1(new_n1052), .B2(new_n829), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1051), .B1(new_n1053), .B2(KEYINPUT50), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT113), .B1(new_n1054), .B2(new_n1048), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT120), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1048), .B1(new_n987), .B2(new_n988), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT120), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n1046), .A4(new_n1049), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1041), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1056), .A2(G168), .A3(new_n1061), .ZN(new_n1063));
  AND2_X1   g638(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1059), .A2(new_n1046), .A3(new_n1049), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(G8), .ZN(new_n1067));
  AOI21_X1  g642(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1062), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT123), .ZN(new_n1074));
  AOI211_X1 g649(.A(new_n1073), .B(G2078), .C1(new_n932), .C2(new_n1074), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n980), .A2(KEYINPUT123), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1075), .A2(new_n977), .A3(new_n1076), .A4(new_n931), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n989), .A2(new_n693), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n1073), .B1(new_n1079), .B2(G2078), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1072), .B1(new_n1081), .B2(G171), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1045), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1073), .A2(G2078), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1083), .A2(new_n980), .A3(new_n1043), .A4(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1078), .A2(KEYINPUT122), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(KEYINPUT122), .B1(new_n1078), .B2(new_n1085), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1080), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1082), .B1(new_n1088), .B2(new_n551), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT124), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  OAI211_X1 g666(.A(KEYINPUT124), .B(new_n1082), .C1(new_n1088), .C2(new_n551), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n977), .A2(new_n980), .A3(new_n978), .ZN(new_n1094));
  OAI22_X1  g669(.A1(new_n989), .A2(G2090), .B1(new_n1094), .B2(G1971), .ZN(new_n1095));
  NAND3_X1  g670(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT55), .ZN(new_n1097));
  INV_X1    g672(.A(G8), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1097), .B1(G166), .B2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1095), .A2(G8), .A3(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1098), .B1(new_n1053), .B2(new_n980), .ZN(new_n1102));
  INV_X1    g677(.A(G1976), .ZN(new_n1103));
  OR2_X1    g678(.A1(G288), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT108), .B(G1976), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT52), .B1(G288), .B2(new_n1105), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1102), .A2(KEYINPUT109), .A3(new_n1104), .A4(new_n1106), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1104), .A2(new_n985), .A3(new_n1106), .A4(G8), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT109), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(G86), .ZN(new_n1111));
  INV_X1    g686(.A(G48), .ZN(new_n1112));
  OAI22_X1  g687(.A1(new_n506), .A2(new_n1111), .B1(new_n508), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n568), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT72), .ZN(new_n1115));
  XNOR2_X1  g690(.A(new_n565), .B(new_n1115), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n495), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(G1981), .B1(new_n1113), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(G1981), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n562), .A2(new_n564), .A3(new_n569), .A4(new_n1119), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1118), .A2(KEYINPUT49), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT49), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1107), .A2(new_n1110), .B1(new_n1102), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1104), .A2(new_n985), .A3(G8), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT52), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1126), .A2(KEYINPUT107), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT107), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1125), .A2(new_n1128), .A3(KEYINPUT52), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n1101), .A2(new_n1124), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1100), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1094), .A2(G1971), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n970), .A2(new_n973), .ZN(new_n1134));
  AOI21_X1  g709(.A(G2090), .B1(new_n1134), .B2(KEYINPUT111), .ZN(new_n1135));
  OR3_X1    g710(.A1(new_n1000), .A2(new_n1001), .A3(KEYINPUT111), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1132), .B1(new_n1137), .B2(new_n1098), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1131), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1088), .A2(new_n551), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1081), .A2(new_n551), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  XOR2_X1   g717(.A(KEYINPUT121), .B(KEYINPUT54), .Z(new_n1143));
  AOI21_X1  g718(.A(new_n1139), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1040), .A2(new_n1071), .A3(new_n1093), .A4(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT125), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1146), .B1(new_n1070), .B2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1131), .A2(new_n1138), .A3(new_n551), .A4(new_n1088), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1149), .B1(new_n1070), .B2(new_n1147), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1063), .A2(new_n1064), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1151));
  OAI211_X1 g726(.A(KEYINPUT125), .B(KEYINPUT62), .C1(new_n1151), .C2(new_n1062), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1148), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1120), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1123), .A2(new_n1102), .ZN(new_n1155));
  NOR2_X1   g730(.A1(G288), .A2(G1976), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT110), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1102), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1161));
  OAI22_X1  g736(.A1(new_n1159), .A2(new_n1160), .B1(new_n1101), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT63), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1066), .A2(G8), .A3(G168), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1163), .B1(new_n1139), .B2(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n1164), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1095), .A2(G8), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1163), .B1(new_n1167), .B2(new_n1132), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1131), .A2(new_n1166), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g744(.A(new_n1162), .B1(new_n1165), .B2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1145), .A2(new_n1153), .A3(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g746(.A(new_n576), .B(new_n948), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n947), .B1(new_n933), .B2(new_n1172), .ZN(new_n1173));
  AND3_X1   g748(.A1(new_n1171), .A2(KEYINPUT126), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT126), .B1(new_n1171), .B2(new_n1173), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n956), .B1(new_n1174), .B2(new_n1175), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g751(.A1(new_n924), .A2(new_n925), .ZN(new_n1178));
  NOR4_X1   g752(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1179));
  OAI21_X1  g753(.A(new_n1179), .B1(new_n853), .B2(new_n854), .ZN(new_n1180));
  NOR2_X1   g754(.A1(new_n1178), .A2(new_n1180), .ZN(G308));
  OAI221_X1 g755(.A(new_n1179), .B1(new_n854), .B2(new_n853), .C1(new_n924), .C2(new_n925), .ZN(G225));
endmodule


