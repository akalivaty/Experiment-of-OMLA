//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:27 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1025, new_n1026, new_n1027, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1048, new_n1049;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n202));
  XNOR2_X1  g001(.A(G8gat), .B(G36gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(G64gat), .ZN(new_n204));
  INV_X1    g003(.A(G92gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(G169gat), .A2(G176gat), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT26), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AND2_X1   g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT27), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT27), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G183gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT28), .ZN(new_n218));
  INV_X1    g017(.A(G190gat), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n215), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n213), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT27), .B(G183gat), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n218), .B1(new_n222), .B2(new_n219), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n214), .A2(new_n219), .ZN(new_n224));
  NOR3_X1   g023(.A1(new_n221), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT25), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n227), .A2(G183gat), .A3(G190gat), .ZN(new_n228));
  XNOR2_X1  g027(.A(G183gat), .B(G190gat), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n228), .B1(new_n229), .B2(new_n227), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n226), .B1(new_n230), .B2(KEYINPUT65), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT64), .B1(new_n207), .B2(KEYINPUT23), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  OAI211_X1 g033(.A(new_n233), .B(new_n234), .C1(G169gat), .C2(G176gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g035(.A1(new_n219), .A2(G183gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n214), .A2(G190gat), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT24), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n210), .B1(KEYINPUT23), .B2(new_n207), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n239), .A2(new_n228), .A3(new_n240), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n231), .A2(new_n236), .A3(new_n241), .ZN(new_n242));
  NAND4_X1  g041(.A1(new_n236), .A2(new_n239), .A3(new_n228), .A4(new_n240), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT65), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n239), .A2(new_n244), .A3(new_n228), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n226), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n225), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G226gat), .ZN(new_n248));
  INV_X1    g047(.A(G233gat), .ZN(new_n249));
  OAI22_X1  g048(.A1(new_n247), .A2(KEYINPUT29), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n242), .A2(new_n246), .ZN(new_n251));
  INV_X1    g050(.A(new_n225), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n248), .A2(new_n249), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G197gat), .B(G204gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT69), .B(G218gat), .ZN(new_n258));
  INV_X1    g057(.A(G211gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n257), .B1(new_n260), .B2(KEYINPUT22), .ZN(new_n261));
  XNOR2_X1  g060(.A(G211gat), .B(G218gat), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(KEYINPUT70), .ZN(new_n263));
  OR2_X1    g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n263), .ZN(new_n265));
  AND2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n256), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n264), .A2(new_n265), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n255), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n206), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT30), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n267), .A2(new_n269), .A3(new_n206), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND4_X1  g072(.A1(new_n267), .A2(KEYINPUT30), .A3(new_n269), .A4(new_n206), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n202), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n272), .A2(new_n271), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n267), .A2(new_n269), .ZN(new_n277));
  INV_X1    g076(.A(new_n206), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n276), .A2(new_n279), .A3(new_n202), .A4(new_n274), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n275), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT79), .ZN(new_n283));
  NAND2_X1  g082(.A1(G225gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT1), .ZN(new_n285));
  XOR2_X1   g084(.A(G113gat), .B(G120gat), .Z(new_n286));
  XOR2_X1   g085(.A(G127gat), .B(G134gat), .Z(new_n287));
  OAI211_X1 g086(.A(new_n285), .B(new_n286), .C1(new_n287), .C2(KEYINPUT66), .ZN(new_n288));
  INV_X1    g087(.A(G113gat), .ZN(new_n289));
  INV_X1    g088(.A(G120gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G113gat), .A2(G120gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(new_n285), .A3(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G127gat), .B(G134gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n291), .A2(new_n292), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n293), .B(new_n294), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n288), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT71), .B1(G155gat), .B2(G162gat), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G155gat), .A2(G162gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NOR3_X1   g102(.A1(KEYINPUT71), .A2(G155gat), .A3(G162gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G141gat), .B(G148gat), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT72), .B(KEYINPUT2), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n303), .B(new_n305), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n306), .ZN(new_n309));
  OR2_X1    g108(.A1(G155gat), .A2(G162gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n301), .ZN(new_n311));
  INV_X1    g110(.A(G155gat), .ZN(new_n312));
  OR2_X1    g111(.A1(KEYINPUT73), .A2(G162gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(KEYINPUT73), .A2(G162gat), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT2), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n309), .B(new_n311), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n308), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n298), .B1(new_n318), .B2(KEYINPUT3), .ZN(new_n319));
  XOR2_X1   g118(.A(KEYINPUT73), .B(G162gat), .Z(new_n320));
  OAI21_X1  g119(.A(KEYINPUT2), .B1(new_n320), .B2(new_n312), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n306), .B1(new_n301), .B2(new_n310), .ZN(new_n322));
  XOR2_X1   g121(.A(KEYINPUT72), .B(KEYINPUT2), .Z(new_n323));
  NAND2_X1  g122(.A1(new_n309), .A2(new_n323), .ZN(new_n324));
  NOR3_X1   g123(.A1(new_n300), .A2(new_n304), .A3(new_n302), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n321), .A2(new_n322), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT3), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n298), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT4), .ZN(new_n330));
  AOI22_X1  g129(.A1(new_n319), .A2(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n288), .A2(new_n297), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT74), .B1(new_n332), .B2(new_n318), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n326), .A2(new_n334), .A3(new_n298), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(KEYINPUT4), .A3(new_n335), .ZN(new_n336));
  AOI211_X1 g135(.A(KEYINPUT39), .B(new_n284), .C1(new_n331), .C2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G57gat), .B(G85gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(G1gat), .B(G29gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n338), .B(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(KEYINPUT75), .B(KEYINPUT0), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n283), .B1(new_n337), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n284), .B1(new_n331), .B2(new_n336), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT39), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n347), .A2(KEYINPUT79), .A3(new_n342), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n335), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n318), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n284), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n352), .A2(KEYINPUT39), .ZN(new_n353));
  OR2_X1    g152(.A1(new_n353), .A2(new_n345), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT40), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n284), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n358), .A2(KEYINPUT5), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n331), .A2(new_n336), .A3(new_n359), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n333), .A2(new_n335), .B1(KEYINPUT4), .B2(new_n284), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n326), .A2(KEYINPUT4), .A3(new_n298), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n332), .B1(new_n326), .B2(new_n327), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n318), .A2(KEYINPUT3), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(KEYINPUT5), .B1(new_n361), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n284), .B1(new_n350), .B2(new_n351), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n360), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n343), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n349), .A2(KEYINPUT40), .A3(new_n354), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n357), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT80), .B1(new_n282), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n266), .B1(KEYINPUT29), .B2(new_n364), .ZN(new_n373));
  NAND2_X1  g172(.A1(G228gat), .A2(G233gat), .ZN(new_n374));
  OR2_X1    g173(.A1(new_n261), .A2(new_n262), .ZN(new_n375));
  AOI21_X1  g174(.A(KEYINPUT29), .B1(new_n261), .B2(new_n262), .ZN(new_n376));
  AOI21_X1  g175(.A(KEYINPUT3), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n373), .B(new_n374), .C1(new_n326), .C2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G78gat), .B(G106gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(new_n379), .B(KEYINPUT31), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT29), .B1(new_n264), .B2(new_n265), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n318), .B1(new_n382), .B2(KEYINPUT3), .ZN(new_n383));
  AND2_X1   g182(.A1(new_n383), .A2(new_n373), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n378), .B(new_n381), .C1(new_n384), .C2(new_n374), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n268), .B1(new_n386), .B2(new_n328), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n377), .A2(new_n326), .ZN(new_n388));
  INV_X1    g187(.A(new_n374), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n387), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n374), .B1(new_n383), .B2(new_n373), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n380), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g191(.A(G22gat), .B(G50gat), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n385), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n393), .B1(new_n385), .B2(new_n392), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT81), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n267), .A2(new_n398), .A3(new_n269), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n250), .A2(new_n255), .A3(KEYINPUT81), .A4(new_n268), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n400), .A2(KEYINPUT37), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT38), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n250), .A2(new_n255), .A3(new_n268), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n268), .B1(new_n250), .B2(new_n255), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT37), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n206), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n402), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT82), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n402), .A2(KEYINPUT82), .A3(new_n407), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n342), .B(new_n360), .C1(new_n366), .C2(new_n367), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n369), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n414), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n332), .A2(new_n318), .A3(KEYINPUT74), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n334), .B1(new_n326), .B2(new_n298), .ZN(new_n418));
  OAI22_X1  g217(.A1(new_n417), .A2(new_n418), .B1(new_n330), .B2(new_n358), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n332), .A2(new_n318), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n328), .A2(new_n319), .B1(new_n420), .B2(KEYINPUT4), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n351), .B1(new_n417), .B2(new_n418), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n358), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n422), .A2(new_n424), .A3(KEYINPUT5), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n342), .B1(new_n425), .B2(new_n360), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n416), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n415), .A2(new_n427), .A3(new_n272), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT38), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n277), .A2(KEYINPUT37), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n407), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n428), .A2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n397), .B1(new_n412), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n276), .A2(new_n274), .A3(new_n279), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(KEYINPUT78), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n280), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT80), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n370), .A2(new_n369), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n357), .A4(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n372), .A2(new_n433), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n416), .A2(new_n426), .ZN(new_n441));
  AOI211_X1 g240(.A(new_n342), .B(new_n414), .C1(new_n425), .C2(new_n360), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT77), .B1(new_n443), .B2(new_n434), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n415), .A2(new_n427), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT77), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n445), .A2(new_n446), .A3(new_n274), .A4(new_n273), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n444), .A2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT36), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n450));
  XOR2_X1   g249(.A(G71gat), .B(G99gat), .Z(new_n451));
  XNOR2_X1  g250(.A(G15gat), .B(G43gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n247), .A2(new_n332), .ZN(new_n454));
  AOI211_X1 g253(.A(new_n298), .B(new_n225), .C1(new_n242), .C2(new_n246), .ZN(new_n455));
  NAND2_X1  g254(.A1(G227gat), .A2(G233gat), .ZN(new_n456));
  NOR3_X1   g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT32), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n453), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n457), .A2(KEYINPUT33), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n450), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n253), .A2(new_n298), .ZN(new_n462));
  INV_X1    g261(.A(new_n456), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n247), .A2(new_n332), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT33), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n465), .A2(KEYINPUT32), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT67), .A4(new_n453), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n453), .A2(KEYINPUT33), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n461), .A2(new_n469), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n462), .A2(new_n464), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT34), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n475), .B1(new_n456), .B2(KEYINPUT68), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n474), .A2(new_n456), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n477), .B1(new_n474), .B2(new_n456), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n473), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(new_n453), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n484), .A2(new_n450), .B1(new_n470), .B2(new_n471), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n481), .B1(new_n485), .B2(new_n469), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n449), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n473), .A2(new_n482), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n485), .A2(new_n469), .A3(new_n481), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT36), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n448), .A2(new_n397), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n396), .A2(new_n488), .A3(new_n489), .ZN(new_n492));
  OAI21_X1  g291(.A(KEYINPUT35), .B1(new_n448), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT35), .ZN(new_n494));
  AND4_X1   g293(.A1(new_n494), .A2(new_n396), .A3(new_n488), .A4(new_n489), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n435), .A2(new_n445), .A3(new_n280), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT83), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n435), .A2(KEYINPUT83), .A3(new_n445), .A4(new_n280), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  AOI22_X1  g299(.A1(new_n440), .A2(new_n491), .B1(new_n493), .B2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n502));
  INV_X1    g301(.A(G22gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G15gat), .ZN(new_n504));
  INV_X1    g303(.A(G15gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G22gat), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(G1gat), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G15gat), .B(G22gat), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n511), .A2(new_n507), .A3(G1gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT16), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n512), .A3(new_n514), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n515), .A2(G8gat), .ZN(new_n516));
  INV_X1    g315(.A(G8gat), .ZN(new_n517));
  AOI22_X1  g316(.A1(new_n508), .A2(new_n509), .B1(new_n511), .B2(new_n513), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n517), .B1(new_n518), .B2(new_n512), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT88), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(G36gat), .ZN(new_n521));
  INV_X1    g320(.A(G29gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT85), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT85), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(G29gat), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n521), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n522), .A2(new_n521), .A3(KEYINPUT14), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT14), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(G29gat), .B2(G36gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g329(.A1(new_n526), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G43gat), .ZN(new_n532));
  INV_X1    g331(.A(G50gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT15), .ZN(new_n535));
  NAND2_X1  g334(.A1(G43gat), .A2(G50gat), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n534), .A2(KEYINPUT86), .A3(new_n535), .A4(new_n536), .ZN(new_n537));
  XNOR2_X1  g336(.A(G43gat), .B(G50gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT84), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n534), .A2(KEYINPUT84), .A3(new_n536), .ZN(new_n541));
  AOI22_X1  g340(.A1(new_n531), .A2(new_n537), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT85), .B(G29gat), .ZN(new_n543));
  OAI211_X1 g342(.A(new_n529), .B(new_n527), .C1(new_n543), .C2(new_n521), .ZN(new_n544));
  AND2_X1   g343(.A1(G43gat), .A2(G50gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(G43gat), .A2(G50gat), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n539), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n547), .A2(new_n541), .A3(KEYINPUT15), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT86), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(new_n538), .B2(KEYINPUT15), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n544), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(KEYINPUT17), .B1(new_n542), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n537), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n548), .B1(new_n544), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n555));
  AND2_X1   g354(.A1(new_n548), .A2(new_n550), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n554), .B(new_n555), .C1(new_n556), .C2(new_n544), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n515), .A2(G8gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT88), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n518), .A2(new_n517), .A3(new_n512), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n520), .A2(new_n552), .A3(new_n557), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G229gat), .A2(G233gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n542), .A2(new_n551), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n558), .A2(new_n560), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n562), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT18), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n558), .B(new_n560), .C1(new_n542), .C2(new_n551), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n566), .A2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n563), .B(KEYINPUT13), .Z(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n562), .A2(KEYINPUT18), .A3(new_n563), .A4(new_n566), .ZN(new_n574));
  XNOR2_X1  g373(.A(G113gat), .B(G141gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT11), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(G169gat), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n575), .A2(KEYINPUT11), .ZN(new_n578));
  INV_X1    g377(.A(G169gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n575), .A2(KEYINPUT11), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(G197gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n577), .A2(new_n581), .A3(G197gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(KEYINPUT12), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT12), .B1(new_n584), .B2(new_n585), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g388(.A1(new_n569), .A2(new_n573), .A3(new_n574), .A4(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n590), .A2(KEYINPUT89), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n574), .A2(new_n573), .ZN(new_n592));
  AOI21_X1  g391(.A(new_n589), .B1(new_n592), .B2(new_n569), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n589), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT89), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n567), .A2(new_n568), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n574), .A2(new_n573), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n595), .B(new_n596), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n502), .B1(new_n594), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n595), .B1(new_n597), .B2(new_n598), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n602), .A2(KEYINPUT89), .A3(new_n590), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n603), .A2(KEYINPUT90), .A3(new_n599), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT94), .B(G183gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G71gat), .B(G78gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(G64gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(G57gat), .ZN(new_n611));
  INV_X1    g410(.A(G57gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(G64gat), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G71gat), .A2(G78gat), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT9), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(KEYINPUT91), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(KEYINPUT92), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n619));
  NOR2_X1   g418(.A1(new_n619), .A2(KEYINPUT91), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n609), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT92), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n623), .B1(new_n611), .B2(new_n613), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n622), .A2(new_n624), .A3(new_n608), .A4(new_n617), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT21), .ZN(new_n627));
  XNOR2_X1  g426(.A(G127gat), .B(G155gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n626), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n629), .B1(new_n626), .B2(new_n627), .ZN(new_n632));
  OAI21_X1  g431(.A(G211gat), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n632), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(new_n259), .A3(new_n630), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n636));
  NAND2_X1  g435(.A1(G231gat), .A2(G233gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  NAND3_X1  g437(.A1(new_n633), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n638), .B1(new_n633), .B2(new_n635), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n621), .A2(KEYINPUT93), .A3(new_n625), .ZN(new_n642));
  AOI21_X1  g441(.A(KEYINPUT93), .B1(new_n621), .B2(new_n625), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n565), .B1(new_n644), .B2(KEYINPUT21), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n640), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n645), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n633), .A2(new_n635), .ZN(new_n648));
  INV_X1    g447(.A(new_n638), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n647), .B1(new_n650), .B2(new_n639), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n607), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n645), .B1(new_n640), .B2(new_n641), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n650), .A2(new_n647), .A3(new_n639), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n653), .A2(new_n654), .A3(new_n606), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(G232gat), .A2(G233gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n657), .B(KEYINPUT95), .Z(new_n658));
  INV_X1    g457(.A(KEYINPUT41), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(G190gat), .B(G218gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  XNOR2_X1  g462(.A(G134gat), .B(G162gat), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT99), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n658), .A2(new_n659), .ZN(new_n667));
  NAND2_X1  g466(.A1(G99gat), .A2(G106gat), .ZN(new_n668));
  INV_X1    g467(.A(G85gat), .ZN(new_n669));
  AOI22_X1  g468(.A1(KEYINPUT8), .A2(new_n668), .B1(new_n669), .B2(new_n205), .ZN(new_n670));
  NAND2_X1  g469(.A1(G85gat), .A2(G92gat), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n671), .A2(KEYINPUT7), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT7), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT96), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT96), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT7), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n671), .B1(new_n674), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT97), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n672), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT96), .B(KEYINPUT7), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n680), .A2(KEYINPUT97), .A3(new_n671), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n670), .B1(new_n679), .B2(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(G99gat), .B(G106gat), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n683), .A2(KEYINPUT98), .ZN(new_n684));
  INV_X1    g483(.A(G99gat), .ZN(new_n685));
  INV_X1    g484(.A(G106gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n687), .A2(new_n688), .A3(new_n668), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n684), .A2(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n682), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(KEYINPUT97), .B1(new_n680), .B2(new_n671), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n674), .A2(new_n676), .ZN(new_n694));
  INV_X1    g493(.A(new_n671), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n678), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n693), .A2(new_n696), .A3(new_n672), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(new_n690), .A3(new_n670), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n667), .B1(new_n699), .B2(new_n564), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n697), .A2(new_n690), .A3(new_n670), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n690), .B1(new_n697), .B2(new_n670), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n703), .A2(new_n552), .A3(new_n557), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n666), .B1(new_n700), .B2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n700), .A2(new_n704), .A3(new_n666), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n665), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n707), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n705), .A3(new_n664), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n663), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n706), .A2(new_n665), .A3(new_n707), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n664), .B1(new_n709), .B2(new_n705), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(new_n713), .A3(new_n662), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n656), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(G230gat), .A2(G233gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT101), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n721));
  OAI21_X1  g520(.A(new_n626), .B1(new_n701), .B2(new_n702), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n621), .A2(new_n625), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n692), .A2(new_n723), .A3(new_n698), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n721), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT93), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n626), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n621), .A2(KEYINPUT93), .A3(new_n625), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n727), .A2(KEYINPUT10), .A3(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n729), .A2(new_n703), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n720), .B1(new_n725), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(KEYINPUT102), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT102), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n733), .B(new_n720), .C1(new_n725), .C2(new_n730), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n722), .A2(new_n724), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n720), .ZN(new_n736));
  XNOR2_X1  g535(.A(G120gat), .B(G148gat), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(G204gat), .ZN(new_n738));
  XNOR2_X1  g537(.A(KEYINPUT103), .B(G176gat), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n738), .B(new_n739), .Z(new_n740));
  NOR2_X1   g539(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n732), .A2(new_n734), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n730), .ZN(new_n743));
  INV_X1    g542(.A(new_n721), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n735), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n719), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n740), .B1(new_n746), .B2(new_n736), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n742), .A2(new_n747), .ZN(new_n748));
  NOR4_X1   g547(.A1(new_n501), .A2(new_n605), .A3(new_n717), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n445), .B(KEYINPUT104), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(KEYINPUT105), .B(G1gat), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1324gat));
  NAND2_X1  g553(.A1(new_n749), .A2(new_n436), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT42), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n513), .A2(new_n517), .ZN(new_n757));
  NOR2_X1   g556(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n758));
  OR2_X1    g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OR3_X1    g558(.A1(new_n755), .A2(new_n756), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n755), .A2(G8gat), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n756), .B1(new_n755), .B2(new_n759), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .ZN(G1325gat));
  NOR2_X1   g562(.A1(new_n483), .A2(new_n486), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n505), .A3(new_n764), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n487), .A2(new_n490), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n749), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n767), .B2(new_n505), .ZN(G1326gat));
  NAND2_X1  g567(.A1(new_n749), .A2(new_n397), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT43), .B(G22gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1327gat));
  NOR2_X1   g570(.A1(new_n501), .A2(new_n605), .ZN(new_n772));
  AND3_X1   g571(.A1(new_n653), .A2(new_n654), .A3(new_n606), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n606), .B1(new_n653), .B2(new_n654), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n748), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(new_n715), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n777), .B(KEYINPUT106), .Z(new_n778));
  NAND2_X1  g577(.A1(new_n772), .A2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n780), .A2(new_n543), .A3(new_n751), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT45), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n603), .A2(new_n599), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n776), .A2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n711), .A2(new_n714), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n440), .A2(new_n491), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n493), .A2(new_n500), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT44), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g591(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n793));
  INV_X1    g592(.A(new_n793), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n501), .A2(new_n787), .A3(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n786), .B1(new_n792), .B2(new_n795), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n796), .A2(new_n750), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n782), .B1(new_n543), .B2(new_n797), .ZN(G1328gat));
  NOR3_X1   g597(.A1(new_n779), .A2(G36gat), .A3(new_n282), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(KEYINPUT46), .ZN(new_n800));
  OAI21_X1  g599(.A(G36gat), .B1(new_n796), .B2(new_n282), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(G1329gat));
  OAI211_X1 g601(.A(new_n766), .B(new_n786), .C1(new_n792), .C2(new_n795), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G43gat), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n780), .A2(new_n532), .A3(new_n764), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT108), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(G1330gat));
  NAND3_X1  g607(.A1(new_n780), .A2(new_n533), .A3(new_n397), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n796), .A2(new_n396), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n809), .B1(new_n810), .B2(new_n533), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT48), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n811), .B(new_n812), .ZN(G1331gat));
  NAND3_X1  g612(.A1(new_n716), .A2(new_n783), .A3(new_n748), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n501), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n751), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g616(.A1(new_n501), .A2(new_n282), .A3(new_n814), .ZN(new_n818));
  NOR2_X1   g617(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n819));
  AND2_X1   g618(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n818), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n821), .B1(new_n818), .B2(new_n819), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n822), .B(KEYINPUT109), .ZN(G1333gat));
  INV_X1    g622(.A(G71gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n815), .A2(new_n824), .A3(new_n764), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n815), .A2(new_n766), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n826), .B2(new_n824), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT110), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT110), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n829), .B(new_n825), .C1(new_n826), .C2(new_n824), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n831), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g631(.A1(new_n815), .A2(new_n397), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g633(.A1(new_n784), .A2(new_n775), .ZN(new_n835));
  AOI21_X1  g634(.A(KEYINPUT51), .B1(new_n790), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n837));
  INV_X1    g636(.A(new_n835), .ZN(new_n838));
  NOR4_X1   g637(.A1(new_n501), .A2(new_n837), .A3(new_n787), .A4(new_n838), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n748), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n751), .A2(new_n669), .ZN(new_n842));
  INV_X1    g641(.A(new_n748), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n838), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n788), .A2(new_n789), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n715), .A3(new_n793), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT44), .B1(new_n501), .B2(new_n787), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n849), .A2(new_n751), .ZN(new_n850));
  OAI22_X1  g649(.A1(new_n841), .A2(new_n842), .B1(new_n850), .B2(new_n669), .ZN(G1336gat));
  NOR2_X1   g650(.A1(new_n282), .A2(G92gat), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n748), .B(new_n852), .C1(new_n836), .C2(new_n839), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n854));
  AOI211_X1 g653(.A(new_n282), .B(new_n845), .C1(new_n847), .C2(new_n848), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n853), .B(new_n854), .C1(new_n855), .C2(new_n205), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT114), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n849), .A2(new_n436), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(G92gat), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n860), .A2(KEYINPUT114), .A3(new_n854), .A4(new_n853), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n282), .A2(G92gat), .A3(new_n843), .ZN(new_n863));
  NOR2_X1   g662(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n865), .B1(new_n790), .B2(new_n835), .ZN(new_n866));
  NOR4_X1   g665(.A1(new_n501), .A2(new_n787), .A3(new_n838), .A4(new_n864), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g669(.A(KEYINPUT113), .B(new_n863), .C1(new_n866), .C2(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT111), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n860), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n859), .A2(KEYINPUT111), .A3(G92gat), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n862), .B1(new_n876), .B2(new_n854), .ZN(G1337gat));
  NAND3_X1  g676(.A1(new_n840), .A2(new_n764), .A3(new_n748), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n766), .A2(G99gat), .ZN(new_n879));
  AOI22_X1  g678(.A1(new_n878), .A2(new_n685), .B1(new_n849), .B2(new_n879), .ZN(G1338gat));
  AOI21_X1  g679(.A(new_n686), .B1(new_n849), .B2(new_n397), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n866), .A2(new_n867), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n396), .A2(G106gat), .A3(new_n843), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n840), .A2(new_n883), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n886), .A2(new_n885), .ZN(new_n887));
  OAI22_X1  g686(.A1(new_n884), .A2(new_n885), .B1(new_n887), .B2(new_n881), .ZN(G1339gat));
  NAND4_X1  g687(.A1(new_n787), .A2(new_n775), .A3(new_n783), .A4(new_n843), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(KEYINPUT115), .ZN(new_n890));
  INV_X1    g689(.A(KEYINPUT115), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n716), .A2(new_n891), .A3(new_n783), .A4(new_n843), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT10), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n642), .A2(new_n643), .A3(new_n895), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n735), .A2(new_n744), .B1(new_n699), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n894), .B1(new_n897), .B2(new_n719), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n732), .A3(new_n734), .ZN(new_n899));
  INV_X1    g698(.A(new_n740), .ZN(new_n900));
  XOR2_X1   g699(.A(KEYINPUT116), .B(KEYINPUT54), .Z(new_n901));
  AOI21_X1  g700(.A(new_n900), .B1(new_n746), .B2(new_n901), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n899), .A2(KEYINPUT55), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n742), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT55), .B1(new_n899), .B2(new_n902), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n584), .A2(new_n585), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n563), .B1(new_n562), .B2(new_n566), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n571), .A2(new_n572), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT117), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT117), .ZN(new_n912));
  OAI211_X1 g711(.A(new_n912), .B(new_n907), .C1(new_n908), .C2(new_n909), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n911), .A2(new_n590), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n906), .A2(new_n715), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n748), .ZN(new_n916));
  INV_X1    g715(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n917), .B1(new_n906), .B2(new_n784), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n915), .B1(new_n918), .B2(new_n715), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n893), .B1(new_n919), .B2(new_n656), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n751), .A2(new_n282), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n764), .A3(new_n396), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n923), .A2(new_n289), .A3(new_n605), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n920), .A2(new_n492), .A3(new_n750), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n925), .A2(new_n282), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n784), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n924), .B1(new_n927), .B2(new_n289), .ZN(G1340gat));
  NOR3_X1   g727(.A1(new_n923), .A2(new_n290), .A3(new_n843), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n926), .A2(new_n748), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n929), .B1(new_n930), .B2(new_n290), .ZN(G1341gat));
  INV_X1    g730(.A(G127gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n926), .A2(new_n932), .A3(new_n775), .ZN(new_n933));
  OAI21_X1  g732(.A(G127gat), .B1(new_n923), .B2(new_n656), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1342gat));
  INV_X1    g734(.A(G134gat), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n282), .A2(new_n715), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT118), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n925), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n939), .A2(KEYINPUT56), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT119), .Z(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(KEYINPUT56), .ZN(new_n942));
  OAI21_X1  g741(.A(G134gat), .B1(new_n923), .B2(new_n787), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(G1343gat));
  NOR2_X1   g743(.A1(new_n766), .A2(new_n396), .ZN(new_n945));
  AND2_X1   g744(.A1(new_n922), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(G141gat), .ZN(new_n947));
  INV_X1    g746(.A(new_n605), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT121), .ZN(new_n951));
  AND3_X1   g750(.A1(new_n603), .A2(KEYINPUT90), .A3(new_n599), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT90), .B1(new_n603), .B2(new_n599), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n952), .A2(new_n953), .A3(new_n904), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n905), .B(new_n955), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n917), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n915), .B1(new_n957), .B2(new_n715), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n893), .B1(new_n958), .B2(new_n656), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT57), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n396), .A2(new_n960), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n951), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n903), .A2(new_n742), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n601), .A2(new_n964), .A3(new_n604), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n905), .A2(new_n955), .ZN(new_n966));
  AOI211_X1 g765(.A(KEYINPUT120), .B(KEYINPUT55), .C1(new_n899), .C2(new_n902), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n916), .B1(new_n965), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(new_n787), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n775), .B1(new_n970), .B2(new_n915), .ZN(new_n971));
  OAI211_X1 g770(.A(KEYINPUT121), .B(new_n961), .C1(new_n971), .C2(new_n893), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n960), .B1(new_n920), .B2(new_n396), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n963), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n921), .A2(new_n766), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(new_n784), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n950), .B1(new_n977), .B2(G141gat), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT58), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT122), .ZN(new_n980));
  AOI21_X1  g779(.A(KEYINPUT58), .B1(new_n949), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n981), .B1(new_n980), .B2(new_n949), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n947), .B1(new_n976), .B2(new_n948), .ZN(new_n983));
  OAI22_X1  g782(.A1(new_n978), .A2(new_n979), .B1(new_n982), .B2(new_n983), .ZN(G1344gat));
  NOR2_X1   g783(.A1(new_n396), .A2(KEYINPUT57), .ZN(new_n985));
  NOR3_X1   g784(.A1(new_n948), .A2(new_n717), .A3(new_n748), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n985), .B1(new_n971), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g786(.A(KEYINPUT57), .B1(new_n920), .B2(new_n396), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n987), .A2(new_n988), .A3(new_n748), .A4(new_n975), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(G148gat), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(KEYINPUT59), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(KEYINPUT124), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT124), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n990), .A2(new_n993), .A3(KEYINPUT59), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n974), .A2(new_n748), .A3(new_n975), .ZN(new_n996));
  INV_X1    g795(.A(G148gat), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n997), .A2(KEYINPUT59), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(KEYINPUT123), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT123), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n996), .A2(new_n1001), .A3(new_n998), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n995), .A2(new_n1000), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n946), .A2(new_n997), .A3(new_n748), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(G1345gat));
  NAND3_X1  g804(.A1(new_n946), .A2(new_n312), .A3(new_n775), .ZN(new_n1006));
  AND2_X1   g805(.A1(new_n976), .A2(new_n775), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1006), .B1(new_n1007), .B2(new_n312), .ZN(G1346gat));
  NOR2_X1   g807(.A1(new_n920), .A2(new_n750), .ZN(new_n1009));
  NAND4_X1  g808(.A1(new_n1009), .A2(new_n320), .A3(new_n938), .A4(new_n945), .ZN(new_n1010));
  AND2_X1   g809(.A1(new_n976), .A2(new_n715), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1010), .B1(new_n1011), .B2(new_n320), .ZN(G1347gat));
  NAND2_X1  g811(.A1(new_n750), .A2(new_n436), .ZN(new_n1013));
  NOR3_X1   g812(.A1(new_n920), .A2(new_n492), .A3(new_n1013), .ZN(new_n1014));
  AOI21_X1  g813(.A(G169gat), .B1(new_n1014), .B2(new_n784), .ZN(new_n1015));
  NOR2_X1   g814(.A1(new_n605), .A2(new_n579), .ZN(new_n1016));
  AOI21_X1  g815(.A(new_n1015), .B1(new_n1014), .B2(new_n1016), .ZN(G1348gat));
  NAND2_X1  g816(.A1(new_n1014), .A2(new_n748), .ZN(new_n1018));
  XNOR2_X1  g817(.A(new_n1018), .B(G176gat), .ZN(G1349gat));
  NAND2_X1  g818(.A1(new_n1014), .A2(new_n775), .ZN(new_n1020));
  OAI22_X1  g819(.A1(new_n1020), .A2(new_n222), .B1(KEYINPUT125), .B2(KEYINPUT60), .ZN(new_n1021));
  AOI21_X1  g820(.A(new_n1021), .B1(new_n214), .B2(new_n1020), .ZN(new_n1022));
  NAND2_X1  g821(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n1023));
  XOR2_X1   g822(.A(new_n1022), .B(new_n1023), .Z(G1350gat));
  NOR2_X1   g823(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n1025));
  AOI21_X1  g824(.A(new_n1025), .B1(new_n1014), .B2(new_n715), .ZN(new_n1026));
  NAND2_X1  g825(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n1027));
  XOR2_X1   g826(.A(new_n1026), .B(new_n1027), .Z(G1351gat));
  NAND2_X1  g827(.A1(new_n987), .A2(new_n988), .ZN(new_n1029));
  NOR3_X1   g828(.A1(new_n1029), .A2(new_n766), .A3(new_n1013), .ZN(new_n1030));
  NAND2_X1  g829(.A1(new_n1030), .A2(new_n948), .ZN(new_n1031));
  AOI21_X1  g830(.A(new_n583), .B1(new_n1031), .B2(KEYINPUT127), .ZN(new_n1032));
  OAI21_X1  g831(.A(new_n1032), .B1(KEYINPUT127), .B2(new_n1031), .ZN(new_n1033));
  NOR4_X1   g832(.A1(new_n920), .A2(new_n396), .A3(new_n766), .A4(new_n1013), .ZN(new_n1034));
  XNOR2_X1  g833(.A(new_n1034), .B(KEYINPUT126), .ZN(new_n1035));
  NAND3_X1  g834(.A1(new_n1035), .A2(new_n583), .A3(new_n784), .ZN(new_n1036));
  NAND2_X1  g835(.A1(new_n1033), .A2(new_n1036), .ZN(G1352gat));
  INV_X1    g836(.A(G204gat), .ZN(new_n1038));
  NAND3_X1  g837(.A1(new_n1034), .A2(new_n1038), .A3(new_n748), .ZN(new_n1039));
  XOR2_X1   g838(.A(new_n1039), .B(KEYINPUT62), .Z(new_n1040));
  NOR4_X1   g839(.A1(new_n1029), .A2(new_n766), .A3(new_n843), .A4(new_n1013), .ZN(new_n1041));
  OAI21_X1  g840(.A(new_n1040), .B1(new_n1038), .B2(new_n1041), .ZN(G1353gat));
  NAND3_X1  g841(.A1(new_n1035), .A2(new_n259), .A3(new_n775), .ZN(new_n1043));
  NAND2_X1  g842(.A1(new_n1030), .A2(new_n775), .ZN(new_n1044));
  AND3_X1   g843(.A1(new_n1044), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1045));
  AOI21_X1  g844(.A(KEYINPUT63), .B1(new_n1044), .B2(G211gat), .ZN(new_n1046));
  OAI21_X1  g845(.A(new_n1043), .B1(new_n1045), .B2(new_n1046), .ZN(G1354gat));
  AOI21_X1  g846(.A(G218gat), .B1(new_n1035), .B2(new_n715), .ZN(new_n1048));
  NOR2_X1   g847(.A1(new_n787), .A2(new_n258), .ZN(new_n1049));
  AOI21_X1  g848(.A(new_n1048), .B1(new_n1030), .B2(new_n1049), .ZN(G1355gat));
endmodule


