//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 1 0 1 0 0 1 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1038,
    new_n1039;
  INV_X1    g000(.A(KEYINPUT100), .ZN(new_n202));
  XNOR2_X1  g001(.A(G43gat), .B(G50gat), .ZN(new_n203));
  AND2_X1   g002(.A1(new_n203), .A2(KEYINPUT15), .ZN(new_n204));
  INV_X1    g003(.A(G43gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G50gat), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT15), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(KEYINPUT96), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT96), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n210));
  AOI22_X1  g009(.A1(KEYINPUT97), .A2(new_n206), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT97), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n203), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G36gat), .ZN(new_n215));
  AND2_X1   g014(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(G29gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n219), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(new_n204), .B1(new_n214), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n204), .A2(new_n221), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT98), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT98), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n211), .A2(new_n213), .B1(new_n218), .B2(new_n220), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n226), .B(new_n223), .C1(new_n227), .C2(new_n204), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT17), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(G8gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(G1gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G1gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT16), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n232), .B1(new_n235), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n238), .ZN(new_n240));
  NOR3_X1   g039(.A1(new_n240), .A2(new_n234), .A3(G8gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT17), .B1(new_n222), .B2(new_n224), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n231), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G229gat), .A2(G233gat), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n242), .B1(new_n225), .B2(new_n228), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(KEYINPUT99), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT99), .ZN(new_n248));
  AOI211_X1 g047(.A(new_n248), .B(new_n242), .C1(new_n225), .C2(new_n228), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n244), .B(new_n245), .C1(new_n247), .C2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT18), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G141gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(G197gat), .ZN(new_n254));
  XOR2_X1   g053(.A(KEYINPUT11), .B(G169gat), .Z(new_n255));
  XNOR2_X1  g054(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(KEYINPUT12), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n246), .B(KEYINPUT99), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n258), .A2(KEYINPUT18), .A3(new_n245), .A4(new_n244), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n225), .A2(new_n242), .A3(new_n228), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n247), .B2(new_n249), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n245), .B(KEYINPUT13), .Z(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n252), .A2(new_n257), .A3(new_n259), .A4(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n250), .A2(new_n251), .B1(new_n261), .B2(new_n262), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n257), .B1(new_n266), .B2(new_n259), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n202), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n252), .A2(new_n259), .A3(new_n263), .ZN(new_n269));
  INV_X1    g068(.A(new_n257), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n271), .A2(KEYINPUT100), .A3(new_n264), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G169gat), .ZN(new_n275));
  INV_X1    g074(.A(G176gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n275), .A2(new_n276), .A3(KEYINPUT71), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT26), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT26), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n279), .A2(new_n275), .A3(new_n276), .A4(KEYINPUT71), .ZN(new_n280));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n278), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(G183gat), .A2(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G190gat), .ZN(new_n285));
  INV_X1    g084(.A(G183gat), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n285), .B1(new_n286), .B2(KEYINPUT27), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT27), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(G183gat), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT28), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT69), .B1(new_n288), .B2(G183gat), .ZN(new_n292));
  AOI21_X1  g091(.A(G190gat), .B1(new_n288), .B2(G183gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n294), .A2(new_n286), .A3(KEYINPUT27), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n292), .A2(new_n293), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n290), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n291), .B1(new_n297), .B2(KEYINPUT70), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT70), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n296), .A2(new_n299), .A3(new_n290), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n284), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n275), .A2(new_n276), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n281), .B1(KEYINPUT66), .B2(KEYINPUT23), .ZN(new_n303));
  NAND2_X1  g102(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n302), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(KEYINPUT65), .A2(G169gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n276), .A2(KEYINPUT23), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n286), .A2(new_n285), .ZN(new_n312));
  NAND3_X1  g111(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n313));
  INV_X1    g112(.A(new_n283), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n312), .B(new_n313), .C1(new_n314), .C2(KEYINPUT24), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n306), .A2(new_n311), .A3(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT25), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n276), .A2(KEYINPUT23), .ZN(new_n318));
  OAI21_X1  g117(.A(KEYINPUT25), .B1(new_n318), .B2(G169gat), .ZN(new_n319));
  OR2_X1    g118(.A1(KEYINPUT66), .A2(KEYINPUT23), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(new_n281), .A3(new_n304), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n319), .B1(new_n302), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(KEYINPUT24), .B1(new_n283), .B2(KEYINPUT67), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT67), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n324), .A2(G183gat), .A3(G190gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n326), .A2(new_n312), .A3(new_n313), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n316), .A2(new_n317), .B1(new_n322), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT76), .B1(new_n301), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n316), .A2(new_n317), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n322), .A2(new_n327), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n296), .A2(new_n299), .A3(new_n290), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n299), .B1(new_n296), .B2(new_n290), .ZN(new_n335));
  NOR3_X1   g134(.A1(new_n334), .A2(new_n335), .A3(new_n291), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n332), .B(new_n333), .C1(new_n336), .C2(new_n284), .ZN(new_n337));
  INV_X1    g136(.A(G226gat), .ZN(new_n338));
  INV_X1    g137(.A(G233gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(KEYINPUT29), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n329), .A2(new_n337), .A3(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT68), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n321), .A2(new_n302), .B1(new_n309), .B2(new_n310), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT25), .B1(new_n344), .B2(new_n315), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n317), .B1(new_n310), .B2(new_n275), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n306), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n312), .A2(new_n313), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n348), .B1(new_n325), .B2(new_n323), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n343), .B1(new_n345), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n330), .A2(KEYINPUT68), .A3(new_n331), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n297), .A2(KEYINPUT70), .ZN(new_n354));
  INV_X1    g153(.A(new_n291), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n354), .A2(new_n300), .A3(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n284), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n353), .A2(new_n340), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G197gat), .B(G204gat), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT22), .ZN(new_n362));
  INV_X1    g161(.A(G211gat), .ZN(new_n363));
  INV_X1    g162(.A(G218gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n362), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(G211gat), .B(G218gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OR2_X1    g168(.A1(new_n369), .A2(KEYINPUT75), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n367), .A2(new_n361), .A3(new_n365), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(KEYINPUT75), .A3(new_n371), .ZN(new_n372));
  AND2_X1   g171(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n360), .A2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n333), .B1(new_n358), .B2(new_n332), .ZN(new_n375));
  NOR3_X1   g174(.A1(new_n301), .A2(KEYINPUT76), .A3(new_n328), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n340), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n370), .A2(new_n372), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n345), .A2(new_n350), .A3(new_n343), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT68), .B1(new_n330), .B2(new_n331), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n358), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n341), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n377), .A2(new_n378), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n374), .A2(new_n383), .A3(KEYINPUT77), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT78), .ZN(new_n385));
  INV_X1    g184(.A(new_n340), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n329), .B2(new_n337), .ZN(new_n387));
  INV_X1    g186(.A(new_n341), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n388), .B1(new_n353), .B2(new_n358), .ZN(new_n389));
  NOR3_X1   g188(.A1(new_n387), .A2(new_n389), .A3(new_n373), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT77), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n384), .A2(new_n385), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n385), .B1(new_n384), .B2(new_n392), .ZN(new_n394));
  OAI21_X1  g193(.A(KEYINPUT37), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT37), .B1(new_n384), .B2(new_n392), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT38), .ZN(new_n397));
  XNOR2_X1  g196(.A(G8gat), .B(G36gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(G64gat), .B(G92gat), .ZN(new_n399));
  XOR2_X1   g198(.A(new_n398), .B(new_n399), .Z(new_n400));
  NOR3_X1   g199(.A1(new_n396), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n395), .A2(new_n401), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n342), .A2(new_n359), .A3(new_n378), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT95), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT95), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n342), .A2(new_n359), .A3(new_n405), .A4(new_n378), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n373), .B1(new_n387), .B2(new_n389), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n404), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT37), .ZN(new_n409));
  INV_X1    g208(.A(new_n400), .ZN(new_n410));
  NOR4_X1   g209(.A1(new_n387), .A2(new_n389), .A3(KEYINPUT77), .A4(new_n373), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n387), .A2(new_n389), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n391), .B1(new_n412), .B2(new_n378), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n411), .B1(new_n413), .B2(new_n374), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n409), .B(new_n410), .C1(new_n414), .C2(KEYINPUT37), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n397), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n402), .A2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G141gat), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT82), .B1(new_n418), .B2(G148gat), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT82), .ZN(new_n420));
  INV_X1    g219(.A(G148gat), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n420), .A2(new_n421), .A3(G141gat), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n419), .B(new_n422), .C1(G141gat), .C2(new_n421), .ZN(new_n423));
  NAND2_X1  g222(.A1(G155gat), .A2(G162gat), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT2), .ZN(new_n425));
  INV_X1    g224(.A(G155gat), .ZN(new_n426));
  INV_X1    g225(.A(G162gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT83), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n428), .A2(new_n429), .A3(new_n424), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n429), .B1(new_n428), .B2(new_n424), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n423), .B(new_n425), .C1(new_n430), .C2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT2), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n418), .A2(G148gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n421), .A2(G141gat), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n428), .A2(KEYINPUT81), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n428), .A2(KEYINPUT81), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n436), .A2(new_n437), .A3(new_n424), .A4(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G120gat), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(G113gat), .ZN(new_n441));
  INV_X1    g240(.A(G113gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(G120gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g243(.A(G127gat), .B(G134gat), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT1), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  XOR2_X1   g246(.A(G127gat), .B(G134gat), .Z(new_n448));
  XNOR2_X1  g247(.A(G113gat), .B(G120gat), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n448), .B1(KEYINPUT1), .B2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n432), .A2(new_n439), .A3(new_n447), .A4(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g252(.A1(new_n432), .A2(new_n439), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n447), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT72), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g256(.A(KEYINPUT72), .B1(new_n450), .B2(new_n447), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n454), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n453), .B1(new_n459), .B2(new_n452), .ZN(new_n460));
  NAND2_X1  g259(.A1(G225gat), .A2(G233gat), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n462), .A2(KEYINPUT5), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT86), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT84), .ZN(new_n465));
  INV_X1    g264(.A(new_n447), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n445), .B1(new_n446), .B2(new_n444), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n465), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n450), .A2(KEYINPUT84), .A3(new_n447), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT3), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(new_n432), .B2(new_n439), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g272(.A(KEYINPUT85), .B(KEYINPUT3), .Z(new_n474));
  NAND3_X1  g273(.A1(new_n432), .A2(new_n439), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n464), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  AND3_X1   g275(.A1(new_n450), .A2(KEYINPUT84), .A3(new_n447), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT84), .B1(new_n450), .B2(new_n447), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n432), .A2(new_n439), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT3), .ZN(new_n481));
  AND4_X1   g280(.A1(new_n464), .A2(new_n479), .A3(new_n481), .A4(new_n475), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n460), .B(new_n463), .C1(new_n476), .C2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G1gat), .B(G29gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT0), .ZN(new_n485));
  XNOR2_X1  g284(.A(G57gat), .B(G85gat), .ZN(new_n486));
  XOR2_X1   g285(.A(new_n485), .B(new_n486), .Z(new_n487));
  OAI211_X1 g286(.A(new_n454), .B(KEYINPUT4), .C1(new_n457), .C2(new_n458), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n462), .B1(new_n451), .B2(new_n452), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n479), .A2(new_n481), .A3(new_n475), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT86), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n464), .A3(new_n475), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n490), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT5), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n451), .B1(new_n470), .B2(new_n454), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n495), .B1(new_n496), .B2(new_n462), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n483), .B(new_n487), .C1(new_n494), .C2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT6), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AND2_X1   g300(.A1(new_n488), .A2(new_n489), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n502), .B1(new_n476), .B2(new_n482), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n497), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n487), .B1(new_n504), .B2(new_n483), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT94), .B1(new_n501), .B2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n483), .B1(new_n494), .B2(new_n498), .ZN(new_n507));
  INV_X1    g306(.A(new_n487), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT94), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n509), .A2(new_n510), .A3(new_n500), .A4(new_n499), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT88), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n513), .B1(new_n505), .B2(KEYINPUT6), .ZN(new_n514));
  AND4_X1   g313(.A1(new_n513), .A2(new_n507), .A3(KEYINPUT6), .A4(new_n508), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n410), .B1(new_n384), .B2(new_n392), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n512), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n417), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT31), .B(G50gat), .ZN(new_n521));
  XNOR2_X1  g320(.A(new_n521), .B(KEYINPUT91), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(G106gat), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G228gat), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n471), .B1(new_n378), .B2(KEYINPUT29), .ZN(new_n526));
  AOI211_X1 g325(.A(new_n525), .B(new_n339), .C1(new_n526), .C2(new_n480), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT29), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n475), .A2(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n373), .B1(KEYINPUT90), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(KEYINPUT90), .B2(new_n529), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n369), .A2(new_n371), .ZN(new_n533));
  AOI21_X1  g332(.A(KEYINPUT89), .B1(new_n533), .B2(new_n528), .ZN(new_n534));
  INV_X1    g333(.A(new_n474), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(KEYINPUT89), .A3(new_n528), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n454), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  AND2_X1   g337(.A1(new_n529), .A2(new_n378), .ZN(new_n539));
  OAI22_X1  g338(.A1(new_n538), .A2(new_n539), .B1(new_n525), .B2(new_n339), .ZN(new_n540));
  INV_X1    g339(.A(G22gat), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n532), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n541), .B1(new_n532), .B2(new_n540), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n543), .A2(new_n544), .A3(G78gat), .ZN(new_n545));
  INV_X1    g344(.A(G78gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n532), .A2(new_n540), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(G22gat), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n546), .B1(new_n548), .B2(new_n542), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n524), .B1(new_n545), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(G78gat), .B1(new_n543), .B2(new_n544), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n548), .A2(new_n546), .A3(new_n542), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n551), .A2(new_n552), .A3(new_n523), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT80), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n517), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n555), .A2(new_n556), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n517), .A2(KEYINPUT80), .A3(KEYINPUT30), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n410), .B1(new_n393), .B2(new_n394), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT79), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n378), .B1(new_n342), .B2(new_n359), .ZN(new_n566));
  NOR3_X1   g365(.A1(new_n390), .A2(new_n391), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(KEYINPUT78), .B1(new_n567), .B2(new_n411), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n384), .A2(new_n385), .A3(new_n392), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT79), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n571), .A3(new_n410), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n563), .B1(new_n565), .B2(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n460), .B1(new_n476), .B2(new_n482), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n462), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n575), .B(KEYINPUT39), .C1(new_n462), .C2(new_n496), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT39), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n574), .A2(new_n577), .A3(new_n462), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n578), .A2(KEYINPUT92), .A3(new_n487), .ZN(new_n579));
  AOI21_X1  g378(.A(KEYINPUT92), .B1(new_n578), .B2(new_n487), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n576), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(KEYINPUT93), .A2(KEYINPUT40), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  OAI221_X1 g382(.A(new_n576), .B1(KEYINPUT93), .B2(KEYINPUT40), .C1(new_n579), .C2(new_n580), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n584), .A3(new_n509), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n520), .B(new_n554), .C1(new_n573), .C2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n587));
  NAND2_X1  g386(.A1(G227gat), .A2(G233gat), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT64), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n457), .A2(new_n458), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n353), .A2(new_n591), .A3(new_n358), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n591), .B1(new_n353), .B2(new_n358), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n590), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n591), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n381), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(new_n589), .A3(new_n592), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(KEYINPUT32), .A3(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT32), .ZN(new_n600));
  OAI211_X1 g399(.A(new_n600), .B(new_n590), .C1(new_n593), .C2(new_n594), .ZN(new_n601));
  AND2_X1   g400(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT33), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G15gat), .B(G43gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT73), .ZN(new_n606));
  INV_X1    g405(.A(G71gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(G99gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n604), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(KEYINPUT74), .B(KEYINPUT34), .Z(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(new_n612), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n604), .A2(new_n614), .A3(new_n610), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n602), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n602), .B1(new_n613), .B2(new_n615), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n587), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n613), .A2(new_n615), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n599), .A2(new_n601), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n622), .A2(KEYINPUT36), .A3(new_n616), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT87), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n501), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n499), .A2(KEYINPUT87), .A3(new_n500), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n509), .A3(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n516), .A2(new_n628), .ZN(new_n629));
  NOR4_X1   g428(.A1(new_n414), .A2(new_n555), .A3(new_n556), .A4(new_n410), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n559), .B1(new_n517), .B2(new_n557), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n571), .B1(new_n570), .B2(new_n410), .ZN(new_n633));
  AOI211_X1 g432(.A(KEYINPUT79), .B(new_n400), .C1(new_n568), .C2(new_n569), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n629), .B(new_n632), .C1(new_n633), .C2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(new_n554), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n624), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n586), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n616), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n554), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT35), .B1(new_n635), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT35), .B1(new_n512), .B2(new_n516), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n573), .A2(new_n554), .A3(new_n639), .A4(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n274), .B1(new_n638), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n629), .ZN(new_n646));
  AND2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT102), .B(G57gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(G64gat), .ZN(new_n649));
  INV_X1    g448(.A(G64gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(G57gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n607), .A2(new_n546), .A3(KEYINPUT9), .ZN(new_n653));
  NAND2_X1  g452(.A1(G71gat), .A2(G78gat), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n657), .A2(new_n607), .A3(new_n546), .ZN(new_n658));
  OAI21_X1  g457(.A(KEYINPUT101), .B1(G71gat), .B2(G78gat), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n658), .A2(new_n654), .A3(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT9), .ZN(new_n661));
  INV_X1    g460(.A(G57gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(G64gat), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n661), .B1(new_n651), .B2(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n656), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT103), .B(KEYINPUT21), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(G231gat), .A2(G233gat), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(new_n671), .B(G127gat), .ZN(new_n672));
  INV_X1    g471(.A(new_n242), .ZN(new_n673));
  INV_X1    g472(.A(new_n667), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n673), .B1(KEYINPUT21), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n672), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g475(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(G155gat), .ZN(new_n678));
  XNOR2_X1  g477(.A(G183gat), .B(G211gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  OR2_X1    g479(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n676), .A2(new_n680), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(G99gat), .A2(G106gat), .ZN(new_n685));
  INV_X1    g484(.A(G85gat), .ZN(new_n686));
  INV_X1    g485(.A(G92gat), .ZN(new_n687));
  AOI22_X1  g486(.A1(KEYINPUT8), .A2(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND3_X1  g489(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n688), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(G106gat), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n609), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n694), .A2(new_n695), .A3(new_n685), .ZN(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n695), .B1(new_n694), .B2(new_n685), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n692), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(G99gat), .B(G106gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(KEYINPUT104), .ZN(new_n701));
  INV_X1    g500(.A(new_n691), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n689), .ZN(new_n703));
  NAND4_X1  g502(.A1(new_n701), .A2(new_n703), .A3(new_n696), .A4(new_n688), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n699), .A2(KEYINPUT105), .A3(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT105), .ZN(new_n706));
  AND4_X1   g505(.A1(new_n701), .A2(new_n703), .A3(new_n696), .A4(new_n688), .ZN(new_n707));
  AOI22_X1  g506(.A1(new_n701), .A2(new_n696), .B1(new_n703), .B2(new_n688), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n706), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n231), .A2(new_n705), .A3(new_n709), .A4(new_n243), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n705), .ZN(new_n711));
  AND2_X1   g510(.A1(G232gat), .A2(G233gat), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n229), .A2(new_n711), .B1(KEYINPUT41), .B2(new_n712), .ZN(new_n713));
  XOR2_X1   g512(.A(G190gat), .B(G218gat), .Z(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n710), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n715), .B1(new_n710), .B2(new_n713), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n712), .A2(KEYINPUT41), .ZN(new_n718));
  XNOR2_X1  g517(.A(G134gat), .B(G162gat), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  OR3_X1    g520(.A1(new_n716), .A2(new_n717), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n716), .B2(new_n717), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(G230gat), .A2(G233gat), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n649), .A2(new_n651), .B1(new_n654), .B2(new_n653), .ZN(new_n727));
  OAI22_X1  g526(.A1(new_n707), .A2(new_n708), .B1(new_n727), .B2(new_n665), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n656), .A2(new_n666), .A3(new_n699), .A4(new_n704), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT10), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n656), .A2(new_n666), .A3(KEYINPUT10), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n731), .B1(new_n709), .B2(new_n705), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n726), .B1(new_n730), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g532(.A(G120gat), .B(G148gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(G176gat), .B(G204gat), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n734), .B(new_n735), .Z(new_n736));
  NAND2_X1  g535(.A1(new_n728), .A2(new_n729), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n733), .B(new_n736), .C1(new_n726), .C2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n737), .A2(new_n726), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n733), .A2(KEYINPUT106), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n741), .B(new_n726), .C1(new_n730), .C2(new_n732), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n739), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n738), .B1(new_n743), .B2(new_n736), .ZN(new_n744));
  NOR3_X1   g543(.A1(new_n684), .A2(new_n725), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n647), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(G1gat), .ZN(G1324gat));
  INV_X1    g546(.A(new_n573), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n645), .A2(new_n745), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G8gat), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT16), .B(G8gat), .Z(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n749), .A2(new_n752), .ZN(new_n753));
  AND3_X1   g552(.A1(new_n753), .A2(KEYINPUT108), .A3(KEYINPUT42), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT108), .B1(new_n753), .B2(KEYINPUT42), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n753), .A2(KEYINPUT42), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n756), .A2(KEYINPUT107), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT107), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n753), .A2(new_n758), .A3(KEYINPUT42), .ZN(new_n759));
  OAI221_X1 g558(.A(new_n750), .B1(new_n754), .B2(new_n755), .C1(new_n757), .C2(new_n759), .ZN(G1325gat));
  AND3_X1   g559(.A1(new_n645), .A2(new_n745), .A3(new_n624), .ZN(new_n761));
  INV_X1    g560(.A(G15gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n645), .A2(new_n639), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n745), .A2(new_n762), .ZN(new_n764));
  OAI22_X1  g563(.A1(new_n761), .A2(new_n762), .B1(new_n763), .B2(new_n764), .ZN(G1326gat));
  NAND3_X1  g564(.A1(new_n645), .A2(new_n745), .A3(new_n636), .ZN(new_n766));
  XNOR2_X1  g565(.A(KEYINPUT43), .B(G22gat), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n766), .B(new_n767), .ZN(G1327gat));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n683), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n681), .A2(KEYINPUT109), .A3(new_n682), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n271), .A2(new_n264), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n773), .A2(new_n744), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n725), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT110), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n635), .A2(new_n636), .ZN(new_n780));
  INV_X1    g579(.A(new_n624), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n565), .A2(new_n572), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n585), .B1(new_n783), .B2(new_n632), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n395), .A2(new_n401), .B1(new_n415), .B2(new_n397), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n512), .A2(new_n516), .A3(new_n518), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n554), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n779), .B1(new_n782), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n586), .A2(new_n637), .A3(KEYINPUT110), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n778), .B1(new_n791), .B2(new_n644), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n638), .A2(new_n644), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n777), .B1(new_n793), .B2(new_n725), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n646), .B(new_n776), .C1(new_n792), .C2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n219), .B1(new_n795), .B2(KEYINPUT111), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n796), .B1(KEYINPUT111), .B2(new_n795), .ZN(new_n797));
  INV_X1    g596(.A(new_n744), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n684), .A2(new_n725), .A3(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n647), .A2(new_n219), .A3(new_n800), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT45), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n797), .A2(new_n802), .ZN(G1328gat));
  OAI211_X1 g602(.A(new_n748), .B(new_n776), .C1(new_n792), .C2(new_n794), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT112), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n215), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n805), .B2(new_n804), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n645), .A2(new_n215), .A3(new_n748), .A4(new_n800), .ZN(new_n808));
  XOR2_X1   g607(.A(new_n808), .B(KEYINPUT46), .Z(new_n809));
  NAND2_X1  g608(.A1(new_n807), .A2(new_n809), .ZN(G1329gat));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n624), .B(new_n776), .C1(new_n792), .C2(new_n794), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n812), .A2(G43gat), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n800), .A2(new_n205), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n763), .A2(new_n814), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n811), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n812), .A2(G43gat), .ZN(new_n817));
  OAI211_X1 g616(.A(new_n817), .B(KEYINPUT47), .C1(new_n763), .C2(new_n814), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(G1330gat));
  NOR2_X1   g618(.A1(new_n799), .A2(G50gat), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n793), .A2(new_n636), .A3(new_n273), .A4(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n636), .B(new_n776), .C1(new_n792), .C2(new_n794), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(G50gat), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT114), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT113), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT48), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AOI211_X1 g628(.A(KEYINPUT114), .B(KEYINPUT48), .C1(new_n821), .C2(new_n826), .ZN(new_n830));
  NOR2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g630(.A(new_n824), .B(new_n831), .ZN(G1331gat));
  AND2_X1   g631(.A1(new_n641), .A2(new_n643), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n833), .B1(new_n789), .B2(new_n790), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n683), .A2(new_n724), .A3(new_n744), .A4(new_n775), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n646), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT115), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n836), .A2(new_n839), .A3(new_n646), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n648), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n841), .B(new_n842), .ZN(G1332gat));
  NAND2_X1  g642(.A1(new_n836), .A2(new_n748), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n844), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT116), .ZN(new_n846));
  XNOR2_X1  g645(.A(KEYINPUT49), .B(G64gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n836), .A2(new_n748), .A3(new_n847), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n845), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n846), .B1(new_n845), .B2(new_n848), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n849), .A2(new_n850), .ZN(G1333gat));
  NAND3_X1  g650(.A1(new_n836), .A2(new_n607), .A3(new_n639), .ZN(new_n852));
  NOR3_X1   g651(.A1(new_n834), .A2(new_n781), .A3(new_n835), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n852), .B1(new_n853), .B2(new_n607), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT50), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n854), .B(new_n855), .ZN(G1334gat));
  NAND2_X1  g655(.A1(new_n836), .A2(new_n636), .ZN(new_n857));
  XNOR2_X1  g656(.A(KEYINPUT117), .B(G78gat), .ZN(new_n858));
  XNOR2_X1  g657(.A(new_n857), .B(new_n858), .ZN(G1335gat));
  NAND2_X1  g658(.A1(new_n684), .A2(new_n775), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT118), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n744), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n586), .A2(new_n637), .A3(KEYINPUT110), .ZN(new_n863));
  AOI21_X1  g662(.A(KEYINPUT110), .B1(new_n586), .B2(new_n637), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n644), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n865), .A2(new_n777), .A3(new_n725), .ZN(new_n866));
  INV_X1    g665(.A(new_n794), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n862), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(G85gat), .B1(new_n869), .B2(new_n629), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n865), .A2(KEYINPUT51), .A3(new_n725), .A4(new_n861), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n861), .A2(new_n725), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n872), .B1(new_n834), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n646), .A2(new_n686), .A3(new_n744), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n870), .B1(new_n876), .B2(new_n877), .ZN(G1336gat));
  INV_X1    g677(.A(KEYINPUT52), .ZN(new_n879));
  INV_X1    g678(.A(new_n862), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n748), .B(new_n880), .C1(new_n792), .C2(new_n794), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n573), .A2(G92gat), .A3(new_n798), .ZN(new_n882));
  XOR2_X1   g681(.A(new_n882), .B(KEYINPUT119), .Z(new_n883));
  AOI22_X1  g682(.A1(new_n881), .A2(G92gat), .B1(new_n875), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n875), .A2(new_n882), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n879), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n687), .B1(new_n868), .B2(new_n748), .ZN(new_n887));
  OAI22_X1  g686(.A1(new_n879), .A2(new_n884), .B1(new_n886), .B2(new_n887), .ZN(G1337gat));
  OAI21_X1  g687(.A(G99gat), .B1(new_n869), .B2(new_n781), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n639), .A2(new_n609), .A3(new_n744), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n876), .B2(new_n890), .ZN(G1338gat));
  AOI21_X1  g690(.A(new_n693), .B1(new_n868), .B2(new_n636), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n636), .A2(new_n693), .A3(new_n744), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n893), .B1(new_n871), .B2(new_n874), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT53), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n636), .B(new_n880), .C1(new_n792), .C2(new_n794), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(G106gat), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT53), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n897), .B(new_n898), .C1(new_n876), .C2(new_n893), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n895), .A2(new_n899), .ZN(G1339gat));
  OR3_X1    g699(.A1(new_n730), .A2(new_n732), .A3(new_n726), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(KEYINPUT54), .A3(new_n733), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n740), .A2(new_n903), .A3(new_n742), .ZN(new_n904));
  INV_X1    g703(.A(new_n736), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n904), .A2(KEYINPUT120), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT120), .B1(new_n904), .B2(new_n905), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT55), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI211_X1 g709(.A(KEYINPUT55), .B(new_n902), .C1(new_n906), .C2(new_n907), .ZN(new_n911));
  NAND4_X1  g710(.A1(new_n910), .A2(new_n774), .A3(new_n738), .A4(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n262), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n258), .A2(new_n260), .A3(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n245), .B1(new_n258), .B2(new_n244), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n256), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n917), .A2(new_n264), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n744), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n725), .B1(new_n912), .B2(new_n919), .ZN(new_n920));
  AND4_X1   g719(.A1(new_n722), .A2(new_n917), .A3(new_n723), .A4(new_n264), .ZN(new_n921));
  AND4_X1   g720(.A1(new_n738), .A2(new_n921), .A3(new_n911), .A4(new_n910), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n772), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n745), .A2(new_n775), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n640), .A2(new_n629), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n573), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n929), .A2(new_n442), .A3(new_n274), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(new_n573), .A3(new_n774), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n930), .B1(new_n442), .B2(new_n931), .ZN(G1340gat));
  NOR2_X1   g731(.A1(new_n929), .A2(new_n798), .ZN(new_n933));
  XNOR2_X1  g732(.A(KEYINPUT121), .B(G120gat), .ZN(new_n934));
  XNOR2_X1  g733(.A(new_n933), .B(new_n934), .ZN(G1341gat));
  OAI21_X1  g734(.A(G127gat), .B1(new_n929), .B2(new_n772), .ZN(new_n936));
  OR2_X1    g735(.A1(new_n684), .A2(G127gat), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n929), .B2(new_n937), .ZN(G1342gat));
  NAND2_X1  g737(.A1(new_n573), .A2(new_n725), .ZN(new_n939));
  NOR3_X1   g738(.A1(new_n927), .A2(G134gat), .A3(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT56), .ZN(new_n941));
  OAI21_X1  g740(.A(G134gat), .B1(new_n929), .B2(new_n724), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1343gat));
  AOI21_X1  g742(.A(new_n554), .B1(new_n923), .B2(new_n924), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT57), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n781), .A2(new_n646), .A3(new_n573), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  AND3_X1   g747(.A1(new_n910), .A2(new_n738), .A3(new_n911), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(new_n921), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n918), .A2(new_n744), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n951), .B1(new_n949), .B2(new_n273), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n950), .B1(new_n952), .B2(new_n725), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n684), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n554), .B1(new_n954), .B2(new_n924), .ZN(new_n955));
  OAI211_X1 g754(.A(new_n946), .B(new_n948), .C1(new_n955), .C2(new_n945), .ZN(new_n956));
  OAI21_X1  g755(.A(G141gat), .B1(new_n956), .B2(new_n274), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT58), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n925), .A2(new_n636), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n959), .A2(new_n947), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n960), .A2(new_n418), .A3(new_n273), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(G141gat), .B1(new_n956), .B2(new_n775), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n963), .A2(new_n961), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n962), .B1(new_n964), .B2(new_n958), .ZN(G1344gat));
  INV_X1    g764(.A(KEYINPUT59), .ZN(new_n966));
  OAI211_X1 g765(.A(new_n966), .B(G148gat), .C1(new_n956), .C2(new_n798), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT123), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n947), .A2(new_n798), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n959), .A2(KEYINPUT57), .ZN(new_n970));
  AND2_X1   g769(.A1(new_n745), .A2(new_n274), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n683), .B1(new_n953), .B2(KEYINPUT122), .ZN(new_n972));
  INV_X1    g771(.A(KEYINPUT122), .ZN(new_n973));
  OAI211_X1 g772(.A(new_n973), .B(new_n950), .C1(new_n952), .C2(new_n725), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n971), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n554), .A2(KEYINPUT57), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n969), .B(new_n970), .C1(new_n975), .C2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(G148gat), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n968), .B1(new_n979), .B2(KEYINPUT59), .ZN(new_n980));
  AOI211_X1 g779(.A(KEYINPUT123), .B(new_n966), .C1(new_n978), .C2(G148gat), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n967), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n944), .A2(new_n969), .A3(new_n421), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(G1345gat));
  NOR3_X1   g783(.A1(new_n956), .A2(new_n426), .A3(new_n772), .ZN(new_n985));
  AOI21_X1  g784(.A(G155gat), .B1(new_n960), .B2(new_n683), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n985), .A2(new_n986), .ZN(G1346gat));
  OAI21_X1  g786(.A(G162gat), .B1(new_n956), .B2(new_n724), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n781), .A2(new_n427), .A3(new_n646), .ZN(new_n989));
  OR2_X1    g788(.A1(new_n989), .A2(new_n939), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n988), .B1(new_n959), .B2(new_n990), .ZN(G1347gat));
  NOR3_X1   g790(.A1(new_n573), .A2(new_n640), .A3(new_n646), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n925), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g792(.A(G169gat), .B1(new_n993), .B2(new_n274), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT124), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n925), .A2(new_n992), .ZN(new_n996));
  NAND3_X1  g795(.A1(new_n996), .A2(new_n309), .A3(new_n774), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n995), .A2(new_n997), .ZN(G1348gat));
  NOR2_X1   g797(.A1(new_n993), .A2(new_n798), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(new_n276), .ZN(G1349gat));
  AOI21_X1  g799(.A(new_n286), .B1(new_n996), .B2(new_n773), .ZN(new_n1001));
  NOR2_X1   g800(.A1(new_n286), .A2(KEYINPUT27), .ZN(new_n1002));
  NOR3_X1   g801(.A1(new_n684), .A2(new_n289), .A3(new_n1002), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n1001), .B1(new_n996), .B2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g803(.A(new_n1004), .B(KEYINPUT60), .Z(G1350gat));
  NAND2_X1  g804(.A1(new_n996), .A2(new_n725), .ZN(new_n1006));
  INV_X1    g805(.A(KEYINPUT125), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n1006), .A2(new_n1007), .A3(G190gat), .ZN(new_n1008));
  NOR2_X1   g807(.A1(new_n993), .A2(new_n724), .ZN(new_n1009));
  OAI21_X1  g808(.A(KEYINPUT125), .B1(new_n1009), .B2(new_n285), .ZN(new_n1010));
  AND3_X1   g809(.A1(new_n1008), .A2(new_n1010), .A3(KEYINPUT61), .ZN(new_n1011));
  OAI22_X1  g810(.A1(new_n1010), .A2(KEYINPUT61), .B1(G190gat), .B2(new_n1006), .ZN(new_n1012));
  OR3_X1    g811(.A1(new_n1011), .A2(new_n1012), .A3(KEYINPUT126), .ZN(new_n1013));
  OAI21_X1  g812(.A(KEYINPUT126), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1013), .A2(new_n1014), .ZN(G1351gat));
  NOR3_X1   g814(.A1(new_n573), .A2(new_n624), .A3(new_n646), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n944), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g816(.A(new_n1017), .ZN(new_n1018));
  AOI21_X1  g817(.A(G197gat), .B1(new_n1018), .B2(new_n774), .ZN(new_n1019));
  NOR2_X1   g818(.A1(new_n975), .A2(new_n977), .ZN(new_n1020));
  INV_X1    g819(.A(new_n970), .ZN(new_n1021));
  INV_X1    g820(.A(new_n1016), .ZN(new_n1022));
  NOR3_X1   g821(.A1(new_n1020), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  AND2_X1   g822(.A1(new_n273), .A2(G197gat), .ZN(new_n1024));
  AOI21_X1  g823(.A(new_n1019), .B1(new_n1023), .B2(new_n1024), .ZN(G1352gat));
  NOR3_X1   g824(.A1(new_n1017), .A2(G204gat), .A3(new_n798), .ZN(new_n1026));
  XNOR2_X1  g825(.A(new_n1026), .B(KEYINPUT62), .ZN(new_n1027));
  NOR4_X1   g826(.A1(new_n1020), .A2(new_n1021), .A3(new_n798), .A4(new_n1022), .ZN(new_n1028));
  AND2_X1   g827(.A1(new_n1028), .A2(KEYINPUT127), .ZN(new_n1029));
  OAI21_X1  g828(.A(G204gat), .B1(new_n1028), .B2(KEYINPUT127), .ZN(new_n1030));
  OAI21_X1  g829(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(G1353gat));
  NAND3_X1  g830(.A1(new_n1018), .A2(new_n363), .A3(new_n683), .ZN(new_n1032));
  INV_X1    g831(.A(new_n1020), .ZN(new_n1033));
  NAND4_X1  g832(.A1(new_n1033), .A2(new_n683), .A3(new_n970), .A4(new_n1016), .ZN(new_n1034));
  AND3_X1   g833(.A1(new_n1034), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1035));
  AOI21_X1  g834(.A(KEYINPUT63), .B1(new_n1034), .B2(G211gat), .ZN(new_n1036));
  OAI21_X1  g835(.A(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(G1354gat));
  NAND3_X1  g836(.A1(new_n1018), .A2(new_n364), .A3(new_n725), .ZN(new_n1038));
  AND2_X1   g837(.A1(new_n1023), .A2(new_n725), .ZN(new_n1039));
  OAI21_X1  g838(.A(new_n1038), .B1(new_n1039), .B2(new_n364), .ZN(G1355gat));
endmodule


