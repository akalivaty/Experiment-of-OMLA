

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U553 ( .A(KEYINPUT102), .ZN(n697) );
  NOR2_X1 U554 ( .A1(G651), .A2(n636), .ZN(n646) );
  AND2_X1 U555 ( .A1(n887), .A2(G126), .ZN(n522) );
  NOR2_X1 U556 ( .A1(n924), .A2(n691), .ZN(n699) );
  INV_X1 U557 ( .A(KEYINPUT29), .ZN(n714) );
  INV_X1 U558 ( .A(KEYINPUT107), .ZN(n732) );
  XNOR2_X1 U559 ( .A(n733), .B(n732), .ZN(n739) );
  XNOR2_X1 U560 ( .A(n539), .B(n538), .ZN(n606) );
  XOR2_X1 U561 ( .A(KEYINPUT1), .B(n523), .Z(n655) );
  AND2_X1 U562 ( .A1(n547), .A2(n546), .ZN(G164) );
  INV_X1 U563 ( .A(G651), .ZN(n527) );
  NOR2_X1 U564 ( .A1(G543), .A2(n527), .ZN(n523) );
  NAND2_X1 U565 ( .A1(G63), .A2(n655), .ZN(n525) );
  XOR2_X1 U566 ( .A(KEYINPUT0), .B(G543), .Z(n636) );
  NAND2_X1 U567 ( .A1(G51), .A2(n646), .ZN(n524) );
  NAND2_X1 U568 ( .A1(n525), .A2(n524), .ZN(n526) );
  XOR2_X1 U569 ( .A(KEYINPUT6), .B(n526), .Z(n535) );
  NOR2_X1 U570 ( .A1(n636), .A2(n527), .ZN(n648) );
  NAND2_X1 U571 ( .A1(G76), .A2(n648), .ZN(n531) );
  XOR2_X1 U572 ( .A(KEYINPUT4), .B(KEYINPUT73), .Z(n529) );
  NOR2_X1 U573 ( .A1(G651), .A2(G543), .ZN(n649) );
  NAND2_X1 U574 ( .A1(G89), .A2(n649), .ZN(n528) );
  XNOR2_X1 U575 ( .A(n529), .B(n528), .ZN(n530) );
  NAND2_X1 U576 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U577 ( .A(n532), .B(KEYINPUT74), .ZN(n533) );
  XNOR2_X1 U578 ( .A(KEYINPUT5), .B(n533), .ZN(n534) );
  NAND2_X1 U579 ( .A1(n535), .A2(n534), .ZN(n536) );
  XNOR2_X1 U580 ( .A(KEYINPUT7), .B(n536), .ZN(G168) );
  XOR2_X1 U581 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  AND2_X1 U582 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U583 ( .A(G57), .ZN(G237) );
  INV_X1 U584 ( .A(G69), .ZN(G235) );
  INV_X1 U585 ( .A(G108), .ZN(G238) );
  INV_X1 U586 ( .A(G120), .ZN(G236) );
  INV_X1 U587 ( .A(G132), .ZN(G219) );
  INV_X1 U588 ( .A(G82), .ZN(G220) );
  NOR2_X1 U589 ( .A1(G2104), .A2(G2105), .ZN(n537) );
  XNOR2_X1 U590 ( .A(n537), .B(KEYINPUT64), .ZN(n539) );
  XNOR2_X1 U591 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n538) );
  NAND2_X1 U592 ( .A1(n606), .A2(G138), .ZN(n541) );
  INV_X1 U593 ( .A(G2105), .ZN(n543) );
  AND2_X1 U594 ( .A1(n543), .A2(G2104), .ZN(n890) );
  NAND2_X1 U595 ( .A1(G102), .A2(n890), .ZN(n540) );
  NAND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U597 ( .A(n542), .B(KEYINPUT88), .Z(n547) );
  NOR2_X1 U598 ( .A1(G2104), .A2(n543), .ZN(n887) );
  AND2_X1 U599 ( .A1(G2104), .A2(G2105), .ZN(n886) );
  NAND2_X1 U600 ( .A1(G114), .A2(n886), .ZN(n544) );
  XNOR2_X1 U601 ( .A(KEYINPUT87), .B(n544), .ZN(n545) );
  NOR2_X1 U602 ( .A1(n522), .A2(n545), .ZN(n546) );
  NAND2_X1 U603 ( .A1(G64), .A2(n655), .ZN(n549) );
  NAND2_X1 U604 ( .A1(G52), .A2(n646), .ZN(n548) );
  NAND2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U606 ( .A(KEYINPUT67), .B(n550), .Z(n555) );
  NAND2_X1 U607 ( .A1(G77), .A2(n648), .ZN(n552) );
  NAND2_X1 U608 ( .A1(G90), .A2(n649), .ZN(n551) );
  NAND2_X1 U609 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U610 ( .A(KEYINPUT9), .B(n553), .Z(n554) );
  NOR2_X1 U611 ( .A1(n555), .A2(n554), .ZN(G171) );
  NAND2_X1 U612 ( .A1(n886), .A2(G113), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G101), .A2(n890), .ZN(n556) );
  XOR2_X1 U614 ( .A(KEYINPUT23), .B(n556), .Z(n557) );
  NAND2_X1 U615 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U616 ( .A1(n887), .A2(G125), .ZN(n560) );
  NAND2_X1 U617 ( .A1(G137), .A2(n606), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n561) );
  NOR2_X1 U619 ( .A1(n562), .A2(n561), .ZN(G160) );
  XOR2_X1 U620 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n564) );
  NAND2_X1 U621 ( .A1(G7), .A2(G661), .ZN(n563) );
  XNOR2_X1 U622 ( .A(n564), .B(n563), .ZN(G223) );
  XOR2_X1 U623 ( .A(G223), .B(KEYINPUT70), .Z(n834) );
  NAND2_X1 U624 ( .A1(n834), .A2(G567), .ZN(n565) );
  XOR2_X1 U625 ( .A(KEYINPUT11), .B(n565), .Z(G234) );
  NAND2_X1 U626 ( .A1(G56), .A2(n655), .ZN(n566) );
  XOR2_X1 U627 ( .A(KEYINPUT14), .B(n566), .Z(n573) );
  NAND2_X1 U628 ( .A1(n648), .A2(G68), .ZN(n567) );
  XNOR2_X1 U629 ( .A(KEYINPUT71), .B(n567), .ZN(n570) );
  NAND2_X1 U630 ( .A1(n649), .A2(G81), .ZN(n568) );
  XOR2_X1 U631 ( .A(KEYINPUT12), .B(n568), .Z(n569) );
  NOR2_X1 U632 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U633 ( .A(n571), .B(KEYINPUT13), .ZN(n572) );
  NOR2_X1 U634 ( .A1(n573), .A2(n572), .ZN(n575) );
  NAND2_X1 U635 ( .A1(n646), .A2(G43), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n575), .A2(n574), .ZN(n924) );
  INV_X1 U637 ( .A(G860), .ZN(n596) );
  OR2_X1 U638 ( .A1(n924), .A2(n596), .ZN(G153) );
  INV_X1 U639 ( .A(G171), .ZN(G301) );
  NAND2_X1 U640 ( .A1(G66), .A2(n655), .ZN(n577) );
  NAND2_X1 U641 ( .A1(G79), .A2(n648), .ZN(n576) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G92), .A2(n649), .ZN(n579) );
  NAND2_X1 U644 ( .A1(G54), .A2(n646), .ZN(n578) );
  NAND2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U647 ( .A(KEYINPUT15), .B(n582), .Z(n583) );
  XNOR2_X2 U648 ( .A(KEYINPUT72), .B(n583), .ZN(n931) );
  INV_X1 U649 ( .A(G868), .ZN(n666) );
  AND2_X1 U650 ( .A1(n931), .A2(n666), .ZN(n585) );
  NOR2_X1 U651 ( .A1(n666), .A2(G301), .ZN(n584) );
  NOR2_X1 U652 ( .A1(n585), .A2(n584), .ZN(G284) );
  NAND2_X1 U653 ( .A1(G78), .A2(n648), .ZN(n587) );
  NAND2_X1 U654 ( .A1(G91), .A2(n649), .ZN(n586) );
  NAND2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n655), .A2(G65), .ZN(n588) );
  XOR2_X1 U657 ( .A(KEYINPUT68), .B(n588), .Z(n589) );
  NOR2_X1 U658 ( .A1(n590), .A2(n589), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n646), .A2(G53), .ZN(n591) );
  NAND2_X1 U660 ( .A1(n592), .A2(n591), .ZN(G299) );
  NOR2_X1 U661 ( .A1(G286), .A2(n666), .ZN(n593) );
  XOR2_X1 U662 ( .A(KEYINPUT75), .B(n593), .Z(n595) );
  NOR2_X1 U663 ( .A1(G868), .A2(G299), .ZN(n594) );
  NOR2_X1 U664 ( .A1(n595), .A2(n594), .ZN(G297) );
  NAND2_X1 U665 ( .A1(n596), .A2(G559), .ZN(n597) );
  NAND2_X1 U666 ( .A1(n597), .A2(n931), .ZN(n598) );
  XNOR2_X1 U667 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U668 ( .A1(G868), .A2(n924), .ZN(n601) );
  NAND2_X1 U669 ( .A1(n931), .A2(G868), .ZN(n599) );
  NOR2_X1 U670 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U671 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U672 ( .A1(G99), .A2(n890), .ZN(n603) );
  NAND2_X1 U673 ( .A1(G111), .A2(n886), .ZN(n602) );
  NAND2_X1 U674 ( .A1(n603), .A2(n602), .ZN(n611) );
  NAND2_X1 U675 ( .A1(G123), .A2(n887), .ZN(n604) );
  XNOR2_X1 U676 ( .A(n604), .B(KEYINPUT18), .ZN(n605) );
  XNOR2_X1 U677 ( .A(n605), .B(KEYINPUT76), .ZN(n608) );
  BUF_X1 U678 ( .A(n606), .Z(n892) );
  NAND2_X1 U679 ( .A1(G135), .A2(n892), .ZN(n607) );
  NAND2_X1 U680 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U681 ( .A(KEYINPUT77), .B(n609), .Z(n610) );
  NOR2_X1 U682 ( .A1(n611), .A2(n610), .ZN(n978) );
  XNOR2_X1 U683 ( .A(n978), .B(G2096), .ZN(n612) );
  XNOR2_X1 U684 ( .A(n612), .B(KEYINPUT78), .ZN(n614) );
  INV_X1 U685 ( .A(G2100), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(G156) );
  NAND2_X1 U687 ( .A1(G559), .A2(n931), .ZN(n664) );
  XNOR2_X1 U688 ( .A(n924), .B(n664), .ZN(n615) );
  NOR2_X1 U689 ( .A1(n615), .A2(G860), .ZN(n623) );
  NAND2_X1 U690 ( .A1(G67), .A2(n655), .ZN(n617) );
  NAND2_X1 U691 ( .A1(G55), .A2(n646), .ZN(n616) );
  NAND2_X1 U692 ( .A1(n617), .A2(n616), .ZN(n622) );
  NAND2_X1 U693 ( .A1(G80), .A2(n648), .ZN(n619) );
  NAND2_X1 U694 ( .A1(G93), .A2(n649), .ZN(n618) );
  NAND2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n620) );
  XOR2_X1 U696 ( .A(KEYINPUT79), .B(n620), .Z(n621) );
  NOR2_X1 U697 ( .A1(n622), .A2(n621), .ZN(n667) );
  XNOR2_X1 U698 ( .A(n623), .B(n667), .ZN(G145) );
  NAND2_X1 U699 ( .A1(n646), .A2(G48), .ZN(n630) );
  NAND2_X1 U700 ( .A1(G61), .A2(n655), .ZN(n625) );
  NAND2_X1 U701 ( .A1(G86), .A2(n649), .ZN(n624) );
  NAND2_X1 U702 ( .A1(n625), .A2(n624), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n648), .A2(G73), .ZN(n626) );
  XOR2_X1 U704 ( .A(KEYINPUT2), .B(n626), .Z(n627) );
  NOR2_X1 U705 ( .A1(n628), .A2(n627), .ZN(n629) );
  NAND2_X1 U706 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U707 ( .A(KEYINPUT81), .B(n631), .Z(G305) );
  NAND2_X1 U708 ( .A1(G49), .A2(n646), .ZN(n633) );
  NAND2_X1 U709 ( .A1(G74), .A2(G651), .ZN(n632) );
  NAND2_X1 U710 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U711 ( .A(KEYINPUT80), .B(n634), .ZN(n635) );
  NOR2_X1 U712 ( .A1(n655), .A2(n635), .ZN(n638) );
  NAND2_X1 U713 ( .A1(n636), .A2(G87), .ZN(n637) );
  NAND2_X1 U714 ( .A1(n638), .A2(n637), .ZN(G288) );
  NAND2_X1 U715 ( .A1(G72), .A2(n648), .ZN(n640) );
  NAND2_X1 U716 ( .A1(G85), .A2(n649), .ZN(n639) );
  NAND2_X1 U717 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U718 ( .A1(G60), .A2(n655), .ZN(n642) );
  NAND2_X1 U719 ( .A1(G47), .A2(n646), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n642), .A2(n641), .ZN(n643) );
  NOR2_X1 U721 ( .A1(n644), .A2(n643), .ZN(n645) );
  XOR2_X1 U722 ( .A(KEYINPUT66), .B(n645), .Z(G290) );
  NAND2_X1 U723 ( .A1(G50), .A2(n646), .ZN(n647) );
  XOR2_X1 U724 ( .A(KEYINPUT82), .B(n647), .Z(n654) );
  NAND2_X1 U725 ( .A1(G75), .A2(n648), .ZN(n651) );
  NAND2_X1 U726 ( .A1(G88), .A2(n649), .ZN(n650) );
  NAND2_X1 U727 ( .A1(n651), .A2(n650), .ZN(n652) );
  XOR2_X1 U728 ( .A(KEYINPUT83), .B(n652), .Z(n653) );
  NOR2_X1 U729 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U730 ( .A1(n655), .A2(G62), .ZN(n656) );
  NAND2_X1 U731 ( .A1(n657), .A2(n656), .ZN(G303) );
  INV_X1 U732 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U733 ( .A(KEYINPUT19), .B(G299), .ZN(n658) );
  XNOR2_X1 U734 ( .A(n658), .B(G305), .ZN(n662) );
  XNOR2_X1 U735 ( .A(G288), .B(n667), .ZN(n660) );
  XNOR2_X1 U736 ( .A(G290), .B(G166), .ZN(n659) );
  XNOR2_X1 U737 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U738 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U739 ( .A(n663), .B(n924), .ZN(n904) );
  XNOR2_X1 U740 ( .A(n664), .B(n904), .ZN(n665) );
  NAND2_X1 U741 ( .A1(n665), .A2(G868), .ZN(n669) );
  NAND2_X1 U742 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U743 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U744 ( .A(KEYINPUT84), .B(n670), .Z(G295) );
  NAND2_X1 U745 ( .A1(G2084), .A2(G2078), .ZN(n671) );
  XNOR2_X1 U746 ( .A(n671), .B(KEYINPUT20), .ZN(n672) );
  XNOR2_X1 U747 ( .A(KEYINPUT85), .B(n672), .ZN(n673) );
  NAND2_X1 U748 ( .A1(n673), .A2(G2090), .ZN(n674) );
  XNOR2_X1 U749 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U750 ( .A1(n675), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U751 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U752 ( .A1(G220), .A2(G219), .ZN(n676) );
  XOR2_X1 U753 ( .A(KEYINPUT22), .B(n676), .Z(n677) );
  NOR2_X1 U754 ( .A1(G218), .A2(n677), .ZN(n678) );
  NAND2_X1 U755 ( .A1(G96), .A2(n678), .ZN(n838) );
  NAND2_X1 U756 ( .A1(n838), .A2(G2106), .ZN(n683) );
  NOR2_X1 U757 ( .A1(G236), .A2(G238), .ZN(n680) );
  NOR2_X1 U758 ( .A1(G235), .A2(G237), .ZN(n679) );
  NAND2_X1 U759 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U760 ( .A(KEYINPUT86), .B(n681), .ZN(n839) );
  NAND2_X1 U761 ( .A1(n839), .A2(G567), .ZN(n682) );
  NAND2_X1 U762 ( .A1(n683), .A2(n682), .ZN(n840) );
  NAND2_X1 U763 ( .A1(G661), .A2(G483), .ZN(n684) );
  NOR2_X1 U764 ( .A1(n840), .A2(n684), .ZN(n837) );
  NAND2_X1 U765 ( .A1(n837), .A2(G36), .ZN(G176) );
  NOR2_X1 U766 ( .A1(G164), .A2(G1384), .ZN(n795) );
  NAND2_X1 U767 ( .A1(G160), .A2(G40), .ZN(n794) );
  INV_X1 U768 ( .A(n794), .ZN(n686) );
  NAND2_X1 U769 ( .A1(n795), .A2(n686), .ZN(n722) );
  XNOR2_X1 U770 ( .A(G1996), .B(KEYINPUT99), .ZN(n950) );
  NOR2_X1 U771 ( .A1(n722), .A2(n950), .ZN(n688) );
  XOR2_X1 U772 ( .A(KEYINPUT26), .B(KEYINPUT100), .Z(n687) );
  XNOR2_X1 U773 ( .A(n688), .B(n687), .ZN(n690) );
  INV_X1 U774 ( .A(n722), .ZN(n716) );
  NAND2_X1 U775 ( .A1(n722), .A2(G1341), .ZN(n689) );
  NAND2_X1 U776 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U777 ( .A1(n699), .A2(n931), .ZN(n692) );
  XOR2_X1 U778 ( .A(KEYINPUT101), .B(n692), .Z(n696) );
  NOR2_X1 U779 ( .A1(n716), .A2(G1348), .ZN(n694) );
  NOR2_X1 U780 ( .A1(G2067), .A2(n722), .ZN(n693) );
  NOR2_X1 U781 ( .A1(n694), .A2(n693), .ZN(n695) );
  NAND2_X1 U782 ( .A1(n696), .A2(n695), .ZN(n698) );
  XNOR2_X1 U783 ( .A(n698), .B(n697), .ZN(n701) );
  NOR2_X1 U784 ( .A1(n699), .A2(n931), .ZN(n700) );
  NOR2_X1 U785 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U786 ( .A(n702), .B(KEYINPUT103), .ZN(n708) );
  NAND2_X1 U787 ( .A1(G2072), .A2(n716), .ZN(n703) );
  XOR2_X1 U788 ( .A(KEYINPUT97), .B(n703), .Z(n704) );
  XNOR2_X1 U789 ( .A(KEYINPUT27), .B(n704), .ZN(n706) );
  XOR2_X1 U790 ( .A(G1956), .B(KEYINPUT98), .Z(n1000) );
  NOR2_X1 U791 ( .A1(n716), .A2(n1000), .ZN(n705) );
  NOR2_X1 U792 ( .A1(n706), .A2(n705), .ZN(n710) );
  INV_X1 U793 ( .A(G299), .ZN(n709) );
  NAND2_X1 U794 ( .A1(n710), .A2(n709), .ZN(n707) );
  NAND2_X1 U795 ( .A1(n708), .A2(n707), .ZN(n713) );
  NOR2_X1 U796 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U797 ( .A(n711), .B(KEYINPUT28), .Z(n712) );
  NAND2_X1 U798 ( .A1(n713), .A2(n712), .ZN(n715) );
  XNOR2_X1 U799 ( .A(n715), .B(n714), .ZN(n720) );
  NAND2_X1 U800 ( .A1(G1961), .A2(n722), .ZN(n718) );
  XOR2_X1 U801 ( .A(G2078), .B(KEYINPUT25), .Z(n953) );
  NAND2_X1 U802 ( .A1(n716), .A2(n953), .ZN(n717) );
  NAND2_X1 U803 ( .A1(n718), .A2(n717), .ZN(n721) );
  OR2_X1 U804 ( .A1(G301), .A2(n721), .ZN(n719) );
  NAND2_X1 U805 ( .A1(n720), .A2(n719), .ZN(n743) );
  NAND2_X1 U806 ( .A1(G301), .A2(n721), .ZN(n728) );
  NAND2_X1 U807 ( .A1(G8), .A2(n722), .ZN(n773) );
  NOR2_X1 U808 ( .A1(G1966), .A2(n773), .ZN(n745) );
  NOR2_X1 U809 ( .A1(G2084), .A2(n722), .ZN(n747) );
  NOR2_X1 U810 ( .A1(n745), .A2(n747), .ZN(n723) );
  NAND2_X1 U811 ( .A1(G8), .A2(n723), .ZN(n724) );
  XNOR2_X1 U812 ( .A(KEYINPUT30), .B(n724), .ZN(n725) );
  NOR2_X1 U813 ( .A1(G168), .A2(n725), .ZN(n726) );
  XOR2_X1 U814 ( .A(KEYINPUT104), .B(n726), .Z(n727) );
  NAND2_X1 U815 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U816 ( .A(n729), .B(KEYINPUT105), .ZN(n730) );
  XOR2_X1 U817 ( .A(KEYINPUT31), .B(n730), .Z(n742) );
  NAND2_X1 U818 ( .A1(n743), .A2(n742), .ZN(n731) );
  NAND2_X1 U819 ( .A1(n731), .A2(G286), .ZN(n733) );
  NOR2_X1 U820 ( .A1(G1971), .A2(n773), .ZN(n734) );
  XNOR2_X1 U821 ( .A(n734), .B(KEYINPUT108), .ZN(n736) );
  NOR2_X1 U822 ( .A1(n722), .A2(G2090), .ZN(n735) );
  NOR2_X1 U823 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U824 ( .A1(G303), .A2(n737), .ZN(n738) );
  NAND2_X1 U825 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U826 ( .A1(n740), .A2(G8), .ZN(n741) );
  XNOR2_X1 U827 ( .A(n741), .B(KEYINPUT32), .ZN(n752) );
  AND2_X1 U828 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U829 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U830 ( .A(KEYINPUT106), .B(n746), .ZN(n750) );
  NAND2_X1 U831 ( .A1(G8), .A2(n747), .ZN(n748) );
  XNOR2_X1 U832 ( .A(KEYINPUT96), .B(n748), .ZN(n749) );
  NAND2_X1 U833 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U834 ( .A1(n752), .A2(n751), .ZN(n759) );
  NOR2_X1 U835 ( .A1(G2090), .A2(G303), .ZN(n753) );
  NAND2_X1 U836 ( .A1(G8), .A2(n753), .ZN(n754) );
  NAND2_X1 U837 ( .A1(n759), .A2(n754), .ZN(n755) );
  NAND2_X1 U838 ( .A1(n755), .A2(n773), .ZN(n770) );
  NOR2_X1 U839 ( .A1(G1976), .A2(G288), .ZN(n762) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n756) );
  NOR2_X1 U841 ( .A1(n762), .A2(n756), .ZN(n943) );
  INV_X1 U842 ( .A(KEYINPUT33), .ZN(n757) );
  AND2_X1 U843 ( .A1(n943), .A2(n757), .ZN(n758) );
  NAND2_X1 U844 ( .A1(n759), .A2(n758), .ZN(n768) );
  NAND2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n932) );
  INV_X1 U846 ( .A(n773), .ZN(n760) );
  AND2_X1 U847 ( .A1(n932), .A2(n760), .ZN(n761) );
  NOR2_X1 U848 ( .A1(KEYINPUT33), .A2(n761), .ZN(n765) );
  NAND2_X1 U849 ( .A1(n762), .A2(KEYINPUT33), .ZN(n763) );
  NOR2_X1 U850 ( .A1(n763), .A2(n773), .ZN(n764) );
  NOR2_X1 U851 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U852 ( .A(G1981), .B(G305), .Z(n925) );
  AND2_X1 U853 ( .A1(n766), .A2(n925), .ZN(n767) );
  NAND2_X1 U854 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U855 ( .A1(n770), .A2(n769), .ZN(n821) );
  NOR2_X1 U856 ( .A1(G1981), .A2(G305), .ZN(n771) );
  XNOR2_X1 U857 ( .A(n771), .B(KEYINPUT24), .ZN(n772) );
  XNOR2_X1 U858 ( .A(n772), .B(KEYINPUT95), .ZN(n774) );
  NOR2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n819) );
  XOR2_X1 U860 ( .A(KEYINPUT38), .B(KEYINPUT93), .Z(n776) );
  NAND2_X1 U861 ( .A1(G105), .A2(n890), .ZN(n775) );
  XNOR2_X1 U862 ( .A(n776), .B(n775), .ZN(n783) );
  NAND2_X1 U863 ( .A1(n886), .A2(G117), .ZN(n778) );
  NAND2_X1 U864 ( .A1(G141), .A2(n892), .ZN(n777) );
  NAND2_X1 U865 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U866 ( .A1(n887), .A2(G129), .ZN(n779) );
  XOR2_X1 U867 ( .A(KEYINPUT92), .B(n779), .Z(n780) );
  NOR2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  NAND2_X1 U869 ( .A1(n783), .A2(n782), .ZN(n883) );
  NOR2_X1 U870 ( .A1(G1996), .A2(n883), .ZN(n975) );
  AND2_X1 U871 ( .A1(n883), .A2(G1996), .ZN(n793) );
  NAND2_X1 U872 ( .A1(G107), .A2(n886), .ZN(n784) );
  XOR2_X1 U873 ( .A(KEYINPUT90), .B(n784), .Z(n789) );
  NAND2_X1 U874 ( .A1(G95), .A2(n890), .ZN(n786) );
  NAND2_X1 U875 ( .A1(G131), .A2(n892), .ZN(n785) );
  NAND2_X1 U876 ( .A1(n786), .A2(n785), .ZN(n787) );
  XOR2_X1 U877 ( .A(KEYINPUT91), .B(n787), .Z(n788) );
  NOR2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n791) );
  NAND2_X1 U879 ( .A1(n887), .A2(G119), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n868) );
  AND2_X1 U881 ( .A1(n868), .A2(G1991), .ZN(n792) );
  NOR2_X1 U882 ( .A1(n793), .A2(n792), .ZN(n984) );
  NOR2_X1 U883 ( .A1(n795), .A2(n794), .ZN(n822) );
  INV_X1 U884 ( .A(n822), .ZN(n796) );
  NOR2_X1 U885 ( .A1(n984), .A2(n796), .ZN(n823) );
  NOR2_X1 U886 ( .A1(G1991), .A2(n868), .ZN(n797) );
  XOR2_X1 U887 ( .A(KEYINPUT109), .B(n797), .Z(n979) );
  NOR2_X1 U888 ( .A1(G1986), .A2(G290), .ZN(n798) );
  NOR2_X1 U889 ( .A1(n979), .A2(n798), .ZN(n799) );
  NOR2_X1 U890 ( .A1(n823), .A2(n799), .ZN(n800) );
  NOR2_X1 U891 ( .A1(n975), .A2(n800), .ZN(n803) );
  XOR2_X1 U892 ( .A(KEYINPUT111), .B(KEYINPUT39), .Z(n801) );
  XNOR2_X1 U893 ( .A(KEYINPUT110), .B(n801), .ZN(n802) );
  XNOR2_X1 U894 ( .A(n803), .B(n802), .ZN(n814) );
  NAND2_X1 U895 ( .A1(G104), .A2(n890), .ZN(n805) );
  NAND2_X1 U896 ( .A1(G140), .A2(n892), .ZN(n804) );
  NAND2_X1 U897 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U898 ( .A(KEYINPUT34), .B(n806), .ZN(n811) );
  NAND2_X1 U899 ( .A1(G116), .A2(n886), .ZN(n808) );
  NAND2_X1 U900 ( .A1(G128), .A2(n887), .ZN(n807) );
  NAND2_X1 U901 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U902 ( .A(KEYINPUT35), .B(n809), .Z(n810) );
  NOR2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n812) );
  XOR2_X1 U904 ( .A(KEYINPUT36), .B(n812), .Z(n869) );
  XOR2_X1 U905 ( .A(G2067), .B(KEYINPUT37), .Z(n815) );
  NAND2_X1 U906 ( .A1(n869), .A2(n815), .ZN(n813) );
  XNOR2_X1 U907 ( .A(n813), .B(KEYINPUT89), .ZN(n982) );
  NAND2_X1 U908 ( .A1(n822), .A2(n982), .ZN(n825) );
  NAND2_X1 U909 ( .A1(n814), .A2(n825), .ZN(n816) );
  OR2_X1 U910 ( .A1(n815), .A2(n869), .ZN(n993) );
  NAND2_X1 U911 ( .A1(n816), .A2(n993), .ZN(n817) );
  NAND2_X1 U912 ( .A1(n817), .A2(n822), .ZN(n830) );
  INV_X1 U913 ( .A(n830), .ZN(n818) );
  OR2_X1 U914 ( .A1(n819), .A2(n818), .ZN(n820) );
  NOR2_X1 U915 ( .A1(n821), .A2(n820), .ZN(n832) );
  XNOR2_X1 U916 ( .A(G1986), .B(G290), .ZN(n937) );
  AND2_X1 U917 ( .A1(n937), .A2(n822), .ZN(n828) );
  INV_X1 U918 ( .A(n823), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U920 ( .A(KEYINPUT94), .B(n826), .ZN(n827) );
  OR2_X1 U921 ( .A1(n828), .A2(n827), .ZN(n829) );
  AND2_X1 U922 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U923 ( .A1(n832), .A2(n831), .ZN(n833) );
  XNOR2_X1 U924 ( .A(n833), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U925 ( .A1(G2106), .A2(n834), .ZN(G217) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U927 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U929 ( .A1(n837), .A2(n836), .ZN(G188) );
  INV_X1 U931 ( .A(G96), .ZN(G221) );
  NOR2_X1 U932 ( .A1(n839), .A2(n838), .ZN(G325) );
  INV_X1 U933 ( .A(G325), .ZN(G261) );
  INV_X1 U934 ( .A(n840), .ZN(G319) );
  XOR2_X1 U935 ( .A(KEYINPUT42), .B(G2072), .Z(n842) );
  XNOR2_X1 U936 ( .A(G2067), .B(G2078), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U938 ( .A(n843), .B(G2100), .Z(n845) );
  XNOR2_X1 U939 ( .A(G2084), .B(G2090), .ZN(n844) );
  XNOR2_X1 U940 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U941 ( .A(G2096), .B(KEYINPUT43), .Z(n847) );
  XNOR2_X1 U942 ( .A(KEYINPUT113), .B(G2678), .ZN(n846) );
  XNOR2_X1 U943 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U944 ( .A(n849), .B(n848), .Z(G227) );
  XNOR2_X1 U945 ( .A(G1981), .B(KEYINPUT114), .ZN(n859) );
  XOR2_X1 U946 ( .A(G1976), .B(G1956), .Z(n851) );
  XNOR2_X1 U947 ( .A(G1966), .B(G1961), .ZN(n850) );
  XNOR2_X1 U948 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U949 ( .A(G1971), .B(G1986), .Z(n853) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1991), .ZN(n852) );
  XNOR2_X1 U951 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U952 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U953 ( .A(G2474), .B(KEYINPUT41), .ZN(n856) );
  XNOR2_X1 U954 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U955 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U956 ( .A1(G124), .A2(n887), .ZN(n860) );
  XNOR2_X1 U957 ( .A(n860), .B(KEYINPUT44), .ZN(n863) );
  NAND2_X1 U958 ( .A1(G112), .A2(n886), .ZN(n861) );
  XOR2_X1 U959 ( .A(KEYINPUT115), .B(n861), .Z(n862) );
  NAND2_X1 U960 ( .A1(n863), .A2(n862), .ZN(n867) );
  NAND2_X1 U961 ( .A1(G100), .A2(n890), .ZN(n865) );
  NAND2_X1 U962 ( .A1(G136), .A2(n892), .ZN(n864) );
  NAND2_X1 U963 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U964 ( .A1(n867), .A2(n866), .ZN(G162) );
  XOR2_X1 U965 ( .A(n869), .B(n868), .Z(n870) );
  XNOR2_X1 U966 ( .A(n870), .B(n978), .ZN(n902) );
  XOR2_X1 U967 ( .A(KEYINPUT48), .B(KEYINPUT119), .Z(n872) );
  XNOR2_X1 U968 ( .A(G160), .B(KEYINPUT46), .ZN(n871) );
  XNOR2_X1 U969 ( .A(n872), .B(n871), .ZN(n873) );
  XOR2_X1 U970 ( .A(n873), .B(G162), .Z(n885) );
  NAND2_X1 U971 ( .A1(G103), .A2(n890), .ZN(n875) );
  NAND2_X1 U972 ( .A1(G139), .A2(n892), .ZN(n874) );
  NAND2_X1 U973 ( .A1(n875), .A2(n874), .ZN(n881) );
  NAND2_X1 U974 ( .A1(n886), .A2(G115), .ZN(n876) );
  XOR2_X1 U975 ( .A(KEYINPUT117), .B(n876), .Z(n878) );
  NAND2_X1 U976 ( .A1(n887), .A2(G127), .ZN(n877) );
  NAND2_X1 U977 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U978 ( .A(KEYINPUT47), .B(n879), .Z(n880) );
  NOR2_X1 U979 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U980 ( .A(KEYINPUT118), .B(n882), .Z(n970) );
  XOR2_X1 U981 ( .A(n883), .B(n970), .Z(n884) );
  XNOR2_X1 U982 ( .A(n885), .B(n884), .ZN(n900) );
  NAND2_X1 U983 ( .A1(G118), .A2(n886), .ZN(n889) );
  NAND2_X1 U984 ( .A1(G130), .A2(n887), .ZN(n888) );
  NAND2_X1 U985 ( .A1(n889), .A2(n888), .ZN(n897) );
  NAND2_X1 U986 ( .A1(n890), .A2(G106), .ZN(n891) );
  XNOR2_X1 U987 ( .A(n891), .B(KEYINPUT116), .ZN(n894) );
  NAND2_X1 U988 ( .A1(G142), .A2(n892), .ZN(n893) );
  NAND2_X1 U989 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U990 ( .A(KEYINPUT45), .B(n895), .Z(n896) );
  NOR2_X1 U991 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U992 ( .A(G164), .B(n898), .Z(n899) );
  XNOR2_X1 U993 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U994 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U995 ( .A1(G37), .A2(n903), .ZN(G395) );
  XNOR2_X1 U996 ( .A(G286), .B(n931), .ZN(n905) );
  XNOR2_X1 U997 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U998 ( .A(n906), .B(G171), .ZN(n907) );
  NOR2_X1 U999 ( .A1(G37), .A2(n907), .ZN(G397) );
  XOR2_X1 U1000 ( .A(KEYINPUT112), .B(G2446), .Z(n909) );
  XNOR2_X1 U1001 ( .A(G2443), .B(G2454), .ZN(n908) );
  XNOR2_X1 U1002 ( .A(n909), .B(n908), .ZN(n910) );
  XOR2_X1 U1003 ( .A(n910), .B(G2451), .Z(n912) );
  XNOR2_X1 U1004 ( .A(G1341), .B(G1348), .ZN(n911) );
  XNOR2_X1 U1005 ( .A(n912), .B(n911), .ZN(n916) );
  XOR2_X1 U1006 ( .A(G2435), .B(G2427), .Z(n914) );
  XNOR2_X1 U1007 ( .A(G2430), .B(G2438), .ZN(n913) );
  XNOR2_X1 U1008 ( .A(n914), .B(n913), .ZN(n915) );
  XOR2_X1 U1009 ( .A(n916), .B(n915), .Z(n917) );
  NAND2_X1 U1010 ( .A1(G14), .A2(n917), .ZN(n923) );
  NAND2_X1 U1011 ( .A1(G319), .A2(n923), .ZN(n920) );
  NOR2_X1 U1012 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1013 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1014 ( .A1(n920), .A2(n919), .ZN(n922) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1016 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1017 ( .A(G225), .ZN(G308) );
  INV_X1 U1018 ( .A(n923), .ZN(G401) );
  XNOR2_X1 U1019 ( .A(G16), .B(KEYINPUT56), .ZN(n948) );
  XNOR2_X1 U1020 ( .A(n924), .B(G1341), .ZN(n930) );
  XNOR2_X1 U1021 ( .A(G1966), .B(G168), .ZN(n926) );
  NAND2_X1 U1022 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1023 ( .A(n927), .B(KEYINPUT125), .ZN(n928) );
  XNOR2_X1 U1024 ( .A(KEYINPUT57), .B(n928), .ZN(n929) );
  NOR2_X1 U1025 ( .A1(n930), .A2(n929), .ZN(n946) );
  XNOR2_X1 U1026 ( .A(n931), .B(G1348), .ZN(n933) );
  NAND2_X1 U1027 ( .A1(n933), .A2(n932), .ZN(n941) );
  XNOR2_X1 U1028 ( .A(G299), .B(G1956), .ZN(n935) );
  AND2_X1 U1029 ( .A1(G1971), .A2(G303), .ZN(n934) );
  NOR2_X1 U1030 ( .A1(n935), .A2(n934), .ZN(n939) );
  XNOR2_X1 U1031 ( .A(G1961), .B(G301), .ZN(n936) );
  NOR2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1034 ( .A1(n941), .A2(n940), .ZN(n942) );
  NAND2_X1 U1035 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1036 ( .A(KEYINPUT126), .B(n944), .Z(n945) );
  NAND2_X1 U1037 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1038 ( .A1(n948), .A2(n947), .ZN(n1028) );
  INV_X1 U1039 ( .A(KEYINPUT55), .ZN(n998) );
  XNOR2_X1 U1040 ( .A(G2090), .B(G35), .ZN(n962) );
  XOR2_X1 U1041 ( .A(G2072), .B(G33), .Z(n949) );
  NAND2_X1 U1042 ( .A1(n949), .A2(G28), .ZN(n959) );
  XNOR2_X1 U1043 ( .A(G32), .B(n950), .ZN(n957) );
  XOR2_X1 U1044 ( .A(G2067), .B(G26), .Z(n952) );
  XOR2_X1 U1045 ( .A(G1991), .B(G25), .Z(n951) );
  NAND2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(G27), .B(n953), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1049 ( .A1(n957), .A2(n956), .ZN(n958) );
  NOR2_X1 U1050 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1051 ( .A(KEYINPUT53), .B(n960), .ZN(n961) );
  NOR2_X1 U1052 ( .A1(n962), .A2(n961), .ZN(n965) );
  XOR2_X1 U1053 ( .A(G2084), .B(G34), .Z(n963) );
  XNOR2_X1 U1054 ( .A(KEYINPUT54), .B(n963), .ZN(n964) );
  NAND2_X1 U1055 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1056 ( .A(n998), .B(n966), .ZN(n968) );
  INV_X1 U1057 ( .A(G29), .ZN(n967) );
  NAND2_X1 U1058 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1059 ( .A1(G11), .A2(n969), .ZN(n1026) );
  XOR2_X1 U1060 ( .A(KEYINPUT52), .B(KEYINPUT124), .Z(n996) );
  XOR2_X1 U1061 ( .A(G164), .B(G2078), .Z(n972) );
  XNOR2_X1 U1062 ( .A(G2072), .B(n970), .ZN(n971) );
  NOR2_X1 U1063 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1064 ( .A(KEYINPUT50), .B(n973), .Z(n992) );
  XOR2_X1 U1065 ( .A(G2090), .B(G162), .Z(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n976) );
  XOR2_X1 U1067 ( .A(KEYINPUT122), .B(n976), .Z(n977) );
  XOR2_X1 U1068 ( .A(KEYINPUT51), .B(n977), .Z(n989) );
  NOR2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1070 ( .A(KEYINPUT120), .B(n980), .Z(n981) );
  NOR2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n986) );
  XOR2_X1 U1073 ( .A(G160), .B(G2084), .Z(n985) );
  NOR2_X1 U1074 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1075 ( .A(KEYINPUT121), .B(n987), .ZN(n988) );
  NOR2_X1 U1076 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(KEYINPUT123), .B(n990), .ZN(n991) );
  NOR2_X1 U1078 ( .A1(n992), .A2(n991), .ZN(n994) );
  NAND2_X1 U1079 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1080 ( .A(n996), .B(n995), .ZN(n997) );
  NAND2_X1 U1081 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1082 ( .A1(n999), .A2(G29), .ZN(n1024) );
  XNOR2_X1 U1083 ( .A(n1000), .B(G20), .ZN(n1004) );
  XNOR2_X1 U1084 ( .A(G1341), .B(G19), .ZN(n1002) );
  XNOR2_X1 U1085 ( .A(G6), .B(G1981), .ZN(n1001) );
  NOR2_X1 U1086 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1087 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XOR2_X1 U1088 ( .A(KEYINPUT59), .B(G1348), .Z(n1005) );
  XNOR2_X1 U1089 ( .A(G4), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1090 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1091 ( .A(KEYINPUT60), .B(n1008), .ZN(n1012) );
  XNOR2_X1 U1092 ( .A(G1966), .B(G21), .ZN(n1010) );
  XNOR2_X1 U1093 ( .A(G1961), .B(G5), .ZN(n1009) );
  NOR2_X1 U1094 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1095 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XNOR2_X1 U1096 ( .A(G1971), .B(G22), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(G23), .B(G1976), .ZN(n1013) );
  NOR2_X1 U1098 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  XOR2_X1 U1099 ( .A(G1986), .B(G24), .Z(n1015) );
  NAND2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(KEYINPUT58), .B(n1017), .ZN(n1018) );
  NOR2_X1 U1102 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1103 ( .A(n1020), .B(KEYINPUT61), .ZN(n1022) );
  XNOR2_X1 U1104 ( .A(G16), .B(KEYINPUT127), .ZN(n1021) );
  NAND2_X1 U1105 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1106 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1107 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1108 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1109 ( .A(KEYINPUT62), .B(n1029), .Z(G311) );
  INV_X1 U1110 ( .A(G311), .ZN(G150) );
endmodule

