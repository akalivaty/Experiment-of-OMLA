

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586;

  XNOR2_X1 U324 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U325 ( .A(n416), .B(KEYINPUT101), .ZN(n417) );
  XOR2_X1 U326 ( .A(n369), .B(n378), .Z(n526) );
  XNOR2_X1 U327 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n469) );
  XNOR2_X1 U328 ( .A(n358), .B(G113GAT), .ZN(n359) );
  XNOR2_X1 U329 ( .A(n470), .B(n469), .ZN(n524) );
  XNOR2_X1 U330 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U331 ( .A(n476), .B(KEYINPUT121), .ZN(n477) );
  XNOR2_X1 U332 ( .A(n408), .B(n407), .ZN(n410) );
  XNOR2_X1 U333 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U334 ( .A(n418), .B(n417), .ZN(n512) );
  XOR2_X1 U335 ( .A(n414), .B(n449), .Z(n555) );
  XNOR2_X1 U336 ( .A(KEYINPUT103), .B(n451), .ZN(n499) );
  XNOR2_X1 U337 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U338 ( .A(n456), .B(G43GAT), .ZN(n457) );
  XNOR2_X1 U339 ( .A(n483), .B(n482), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n458), .B(n457), .ZN(G1330GAT) );
  XOR2_X1 U341 ( .A(G85GAT), .B(G162GAT), .Z(n293) );
  XNOR2_X1 U342 ( .A(G148GAT), .B(G155GAT), .ZN(n292) );
  XNOR2_X1 U343 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U344 ( .A(n294), .B(G127GAT), .Z(n296) );
  XOR2_X1 U345 ( .A(G113GAT), .B(G1GAT), .Z(n443) );
  XNOR2_X1 U346 ( .A(G29GAT), .B(n443), .ZN(n295) );
  XNOR2_X1 U347 ( .A(n296), .B(n295), .ZN(n313) );
  XOR2_X1 U348 ( .A(G134GAT), .B(KEYINPUT76), .Z(n394) );
  XOR2_X1 U349 ( .A(KEYINPUT5), .B(G57GAT), .Z(n298) );
  XNOR2_X1 U350 ( .A(KEYINPUT93), .B(KEYINPUT1), .ZN(n297) );
  XNOR2_X1 U351 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U352 ( .A(KEYINPUT98), .B(KEYINPUT94), .Z(n300) );
  XNOR2_X1 U353 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n299) );
  XNOR2_X1 U354 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U355 ( .A(n302), .B(n301), .Z(n307) );
  XOR2_X1 U356 ( .A(KEYINPUT6), .B(KEYINPUT4), .Z(n304) );
  NAND2_X1 U357 ( .A1(G225GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U359 ( .A(KEYINPUT97), .B(n305), .ZN(n306) );
  XNOR2_X1 U360 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U361 ( .A(n394), .B(n308), .Z(n311) );
  XOR2_X1 U362 ( .A(KEYINPUT0), .B(G120GAT), .Z(n356) );
  XNOR2_X1 U363 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n309) );
  XNOR2_X1 U364 ( .A(n309), .B(KEYINPUT2), .ZN(n342) );
  XNOR2_X1 U365 ( .A(n356), .B(n342), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U367 ( .A(n313), .B(n312), .ZN(n513) );
  INV_X1 U368 ( .A(n513), .ZN(n474) );
  XOR2_X1 U369 ( .A(G15GAT), .B(G127GAT), .Z(n357) );
  XNOR2_X1 U370 ( .A(G1GAT), .B(n357), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n314), .B(G64GAT), .ZN(n329) );
  XNOR2_X1 U372 ( .A(G22GAT), .B(G155GAT), .ZN(n315) );
  XNOR2_X1 U373 ( .A(n315), .B(G78GAT), .ZN(n343) );
  XOR2_X1 U374 ( .A(KEYINPUT81), .B(n343), .Z(n317) );
  NAND2_X1 U375 ( .A1(G231GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U376 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U377 ( .A(KEYINPUT14), .B(KEYINPUT80), .Z(n319) );
  XNOR2_X1 U378 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n318) );
  XNOR2_X1 U379 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U380 ( .A(n321), .B(n320), .Z(n327) );
  XOR2_X1 U381 ( .A(KEYINPUT72), .B(KEYINPUT13), .Z(n323) );
  XNOR2_X1 U382 ( .A(G71GAT), .B(G57GAT), .ZN(n322) );
  XNOR2_X1 U383 ( .A(n323), .B(n322), .ZN(n431) );
  XOR2_X1 U384 ( .A(KEYINPUT79), .B(G211GAT), .Z(n325) );
  XNOR2_X1 U385 ( .A(G8GAT), .B(G183GAT), .ZN(n324) );
  XNOR2_X1 U386 ( .A(n325), .B(n324), .ZN(n372) );
  XNOR2_X1 U387 ( .A(n431), .B(n372), .ZN(n326) );
  XNOR2_X1 U388 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U389 ( .A(n329), .B(n328), .Z(n579) );
  XOR2_X1 U390 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n331) );
  XNOR2_X1 U391 ( .A(G197GAT), .B(G218GAT), .ZN(n330) );
  XNOR2_X1 U392 ( .A(n331), .B(n330), .ZN(n379) );
  XNOR2_X1 U393 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n332), .B(G148GAT), .ZN(n423) );
  XNOR2_X1 U395 ( .A(n379), .B(n423), .ZN(n347) );
  XOR2_X1 U396 ( .A(G50GAT), .B(G162GAT), .Z(n397) );
  XOR2_X1 U397 ( .A(G204GAT), .B(G211GAT), .Z(n334) );
  XNOR2_X1 U398 ( .A(KEYINPUT24), .B(KEYINPUT92), .ZN(n333) );
  XNOR2_X1 U399 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U400 ( .A(n397), .B(n335), .Z(n337) );
  NAND2_X1 U401 ( .A1(G228GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U403 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n339) );
  XNOR2_X1 U404 ( .A(KEYINPUT89), .B(KEYINPUT22), .ZN(n338) );
  XNOR2_X1 U405 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U406 ( .A(n341), .B(n340), .Z(n345) );
  XNOR2_X1 U407 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U408 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U409 ( .A(n347), .B(n346), .ZN(n475) );
  XOR2_X1 U410 ( .A(G176GAT), .B(G183GAT), .Z(n349) );
  XNOR2_X1 U411 ( .A(KEYINPUT20), .B(KEYINPUT83), .ZN(n348) );
  XNOR2_X1 U412 ( .A(n349), .B(n348), .ZN(n364) );
  XOR2_X1 U413 ( .A(G99GAT), .B(G134GAT), .Z(n351) );
  XNOR2_X1 U414 ( .A(G43GAT), .B(G190GAT), .ZN(n350) );
  XNOR2_X1 U415 ( .A(n351), .B(n350), .ZN(n355) );
  XOR2_X1 U416 ( .A(G71GAT), .B(KEYINPUT85), .Z(n353) );
  XNOR2_X1 U417 ( .A(KEYINPUT84), .B(KEYINPUT88), .ZN(n352) );
  XNOR2_X1 U418 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U419 ( .A(n355), .B(n354), .Z(n362) );
  XOR2_X1 U420 ( .A(n357), .B(n356), .Z(n360) );
  NAND2_X1 U421 ( .A1(G227GAT), .A2(G233GAT), .ZN(n358) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n369) );
  XOR2_X1 U424 ( .A(KEYINPUT86), .B(KEYINPUT19), .Z(n366) );
  XNOR2_X1 U425 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n365) );
  XNOR2_X1 U426 ( .A(n366), .B(n365), .ZN(n368) );
  XOR2_X1 U427 ( .A(KEYINPUT87), .B(KEYINPUT17), .Z(n367) );
  XOR2_X1 U428 ( .A(n368), .B(n367), .Z(n378) );
  INV_X1 U429 ( .A(n526), .ZN(n455) );
  NOR2_X1 U430 ( .A1(n475), .A2(n455), .ZN(n370) );
  XNOR2_X1 U431 ( .A(n370), .B(KEYINPUT26), .ZN(n569) );
  XNOR2_X1 U432 ( .A(G36GAT), .B(G190GAT), .ZN(n371) );
  XNOR2_X1 U433 ( .A(n371), .B(KEYINPUT78), .ZN(n405) );
  XOR2_X1 U434 ( .A(n372), .B(n405), .Z(n374) );
  NAND2_X1 U435 ( .A1(G226GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U436 ( .A(n374), .B(n373), .ZN(n377) );
  XOR2_X1 U437 ( .A(G64GAT), .B(G92GAT), .Z(n376) );
  XNOR2_X1 U438 ( .A(G176GAT), .B(G204GAT), .ZN(n375) );
  XNOR2_X1 U439 ( .A(n376), .B(n375), .ZN(n422) );
  XOR2_X1 U440 ( .A(n377), .B(n422), .Z(n382) );
  INV_X1 U441 ( .A(n378), .ZN(n380) );
  XOR2_X1 U442 ( .A(n380), .B(n379), .Z(n381) );
  XOR2_X1 U443 ( .A(n382), .B(n381), .Z(n497) );
  XOR2_X1 U444 ( .A(n497), .B(KEYINPUT99), .Z(n383) );
  XNOR2_X1 U445 ( .A(n383), .B(KEYINPUT27), .ZN(n390) );
  NAND2_X1 U446 ( .A1(n569), .A2(n390), .ZN(n387) );
  NAND2_X1 U447 ( .A1(n455), .A2(n497), .ZN(n384) );
  NAND2_X1 U448 ( .A1(n475), .A2(n384), .ZN(n385) );
  XOR2_X1 U449 ( .A(KEYINPUT25), .B(n385), .Z(n386) );
  NAND2_X1 U450 ( .A1(n387), .A2(n386), .ZN(n388) );
  NAND2_X1 U451 ( .A1(n388), .A2(n513), .ZN(n389) );
  XNOR2_X1 U452 ( .A(n389), .B(KEYINPUT100), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n475), .B(KEYINPUT28), .ZN(n520) );
  INV_X1 U454 ( .A(n520), .ZN(n529) );
  NAND2_X1 U455 ( .A1(n474), .A2(n390), .ZN(n523) );
  NOR2_X1 U456 ( .A1(n529), .A2(n523), .ZN(n391) );
  NAND2_X1 U457 ( .A1(n391), .A2(n526), .ZN(n392) );
  NAND2_X1 U458 ( .A1(n393), .A2(n392), .ZN(n487) );
  XOR2_X1 U459 ( .A(G99GAT), .B(G85GAT), .Z(n426) );
  XNOR2_X1 U460 ( .A(n426), .B(n394), .ZN(n396) );
  AND2_X1 U461 ( .A1(G232GAT), .A2(G233GAT), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n396), .B(n395), .ZN(n398) );
  XNOR2_X1 U463 ( .A(n398), .B(n397), .ZN(n408) );
  XOR2_X1 U464 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n400) );
  XNOR2_X1 U465 ( .A(G218GAT), .B(KEYINPUT77), .ZN(n399) );
  XNOR2_X1 U466 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U467 ( .A(KEYINPUT9), .B(KEYINPUT66), .Z(n402) );
  XNOR2_X1 U468 ( .A(KEYINPUT10), .B(KEYINPUT74), .ZN(n401) );
  XNOR2_X1 U469 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U470 ( .A(n404), .B(n403), .Z(n406) );
  XOR2_X1 U471 ( .A(G106GAT), .B(G92GAT), .Z(n409) );
  XNOR2_X1 U472 ( .A(n410), .B(n409), .ZN(n414) );
  XOR2_X1 U473 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n412) );
  XNOR2_X1 U474 ( .A(G43GAT), .B(G29GAT), .ZN(n411) );
  XNOR2_X1 U475 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U476 ( .A(KEYINPUT7), .B(n413), .ZN(n449) );
  INV_X1 U477 ( .A(n555), .ZN(n484) );
  XOR2_X1 U478 ( .A(n484), .B(KEYINPUT36), .Z(n582) );
  NAND2_X1 U479 ( .A1(n487), .A2(n582), .ZN(n415) );
  NOR2_X1 U480 ( .A1(n579), .A2(n415), .ZN(n418) );
  XNOR2_X1 U481 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n416) );
  XOR2_X1 U482 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n420) );
  NAND2_X1 U483 ( .A1(G230GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U484 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U485 ( .A(n421), .B(KEYINPUT31), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n427), .B(n426), .ZN(n429) );
  XNOR2_X1 U489 ( .A(G120GAT), .B(G78GAT), .ZN(n428) );
  XNOR2_X1 U490 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U491 ( .A(n431), .B(n430), .ZN(n574) );
  XOR2_X1 U492 ( .A(KEYINPUT69), .B(KEYINPUT29), .Z(n433) );
  XNOR2_X1 U493 ( .A(KEYINPUT71), .B(KEYINPUT67), .ZN(n432) );
  XNOR2_X1 U494 ( .A(n433), .B(n432), .ZN(n447) );
  XOR2_X1 U495 ( .A(G15GAT), .B(G50GAT), .Z(n435) );
  XNOR2_X1 U496 ( .A(G169GAT), .B(G36GAT), .ZN(n434) );
  XNOR2_X1 U497 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U498 ( .A(G8GAT), .B(G141GAT), .Z(n437) );
  XNOR2_X1 U499 ( .A(G197GAT), .B(G22GAT), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U501 ( .A(n439), .B(n438), .Z(n445) );
  XOR2_X1 U502 ( .A(KEYINPUT30), .B(KEYINPUT68), .Z(n441) );
  NAND2_X1 U503 ( .A1(G229GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U504 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U505 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n446) );
  XOR2_X1 U507 ( .A(n447), .B(n446), .Z(n448) );
  XOR2_X1 U508 ( .A(n449), .B(n448), .Z(n571) );
  INV_X1 U509 ( .A(n571), .ZN(n558) );
  AND2_X1 U510 ( .A1(n574), .A2(n558), .ZN(n489) );
  NAND2_X1 U511 ( .A1(n512), .A2(n489), .ZN(n450) );
  XNOR2_X1 U512 ( .A(n450), .B(KEYINPUT38), .ZN(n451) );
  NAND2_X1 U513 ( .A1(n474), .A2(n499), .ZN(n454) );
  XOR2_X1 U514 ( .A(KEYINPUT39), .B(KEYINPUT104), .Z(n452) );
  XNOR2_X1 U515 ( .A(n452), .B(G29GAT), .ZN(n453) );
  XNOR2_X1 U516 ( .A(n454), .B(n453), .ZN(G1328GAT) );
  NAND2_X1 U517 ( .A1(n455), .A2(n499), .ZN(n458) );
  XOR2_X1 U518 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n456) );
  INV_X1 U519 ( .A(KEYINPUT54), .ZN(n472) );
  XOR2_X1 U520 ( .A(n574), .B(KEYINPUT41), .Z(n532) );
  NOR2_X1 U521 ( .A1(n571), .A2(n532), .ZN(n459) );
  XNOR2_X1 U522 ( .A(n459), .B(KEYINPUT46), .ZN(n460) );
  XOR2_X1 U523 ( .A(KEYINPUT109), .B(n579), .Z(n564) );
  NOR2_X1 U524 ( .A1(n460), .A2(n564), .ZN(n461) );
  NAND2_X1 U525 ( .A1(n461), .A2(n484), .ZN(n462) );
  XNOR2_X1 U526 ( .A(KEYINPUT47), .B(n462), .ZN(n468) );
  XOR2_X1 U527 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n464) );
  NAND2_X1 U528 ( .A1(n579), .A2(n582), .ZN(n463) );
  XNOR2_X1 U529 ( .A(n464), .B(n463), .ZN(n466) );
  NAND2_X1 U530 ( .A1(n571), .A2(n574), .ZN(n465) );
  NOR2_X1 U531 ( .A1(n466), .A2(n465), .ZN(n467) );
  NOR2_X1 U532 ( .A1(n468), .A2(n467), .ZN(n470) );
  INV_X1 U533 ( .A(n497), .ZN(n515) );
  NOR2_X1 U534 ( .A1(n524), .A2(n515), .ZN(n471) );
  XNOR2_X1 U535 ( .A(n472), .B(n471), .ZN(n473) );
  NOR2_X1 U536 ( .A1(n474), .A2(n473), .ZN(n570) );
  AND2_X1 U537 ( .A1(n570), .A2(n475), .ZN(n478) );
  INV_X1 U538 ( .A(KEYINPUT55), .ZN(n476) );
  NOR2_X1 U539 ( .A1(n526), .A2(n479), .ZN(n565) );
  NAND2_X1 U540 ( .A1(n565), .A2(n555), .ZN(n483) );
  XOR2_X1 U541 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n481) );
  XNOR2_X1 U542 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n480) );
  XOR2_X1 U543 ( .A(KEYINPUT16), .B(KEYINPUT82), .Z(n486) );
  NAND2_X1 U544 ( .A1(n579), .A2(n484), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(n488) );
  AND2_X1 U546 ( .A1(n488), .A2(n487), .ZN(n502) );
  NAND2_X1 U547 ( .A1(n489), .A2(n502), .ZN(n495) );
  NOR2_X1 U548 ( .A1(n513), .A2(n495), .ZN(n490) );
  XOR2_X1 U549 ( .A(G1GAT), .B(n490), .Z(n491) );
  XNOR2_X1 U550 ( .A(KEYINPUT34), .B(n491), .ZN(G1324GAT) );
  NOR2_X1 U551 ( .A1(n515), .A2(n495), .ZN(n492) );
  XOR2_X1 U552 ( .A(G8GAT), .B(n492), .Z(G1325GAT) );
  NOR2_X1 U553 ( .A1(n526), .A2(n495), .ZN(n494) );
  XNOR2_X1 U554 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1326GAT) );
  NOR2_X1 U556 ( .A1(n520), .A2(n495), .ZN(n496) );
  XOR2_X1 U557 ( .A(G22GAT), .B(n496), .Z(G1327GAT) );
  NAND2_X1 U558 ( .A1(n499), .A2(n497), .ZN(n498) );
  XNOR2_X1 U559 ( .A(n498), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U560 ( .A1(n499), .A2(n529), .ZN(n500) );
  XNOR2_X1 U561 ( .A(n500), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U562 ( .A1(n532), .A2(n558), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n501), .B(KEYINPUT106), .ZN(n511) );
  NAND2_X1 U564 ( .A1(n502), .A2(n511), .ZN(n508) );
  NOR2_X1 U565 ( .A1(n513), .A2(n508), .ZN(n503) );
  XOR2_X1 U566 ( .A(G57GAT), .B(n503), .Z(n504) );
  XNOR2_X1 U567 ( .A(KEYINPUT42), .B(n504), .ZN(G1332GAT) );
  NOR2_X1 U568 ( .A1(n515), .A2(n508), .ZN(n506) );
  XNOR2_X1 U569 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(G1333GAT) );
  NOR2_X1 U571 ( .A1(n526), .A2(n508), .ZN(n507) );
  XOR2_X1 U572 ( .A(G71GAT), .B(n507), .Z(G1334GAT) );
  NOR2_X1 U573 ( .A1(n520), .A2(n508), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U575 ( .A(n510), .B(n509), .ZN(G1335GAT) );
  NAND2_X1 U576 ( .A1(n512), .A2(n511), .ZN(n519) );
  NOR2_X1 U577 ( .A1(n513), .A2(n519), .ZN(n514) );
  XOR2_X1 U578 ( .A(G85GAT), .B(n514), .Z(G1336GAT) );
  NOR2_X1 U579 ( .A1(n515), .A2(n519), .ZN(n516) );
  XOR2_X1 U580 ( .A(G92GAT), .B(n516), .Z(G1337GAT) );
  NOR2_X1 U581 ( .A1(n526), .A2(n519), .ZN(n517) );
  XOR2_X1 U582 ( .A(KEYINPUT108), .B(n517), .Z(n518) );
  XNOR2_X1 U583 ( .A(G99GAT), .B(n518), .ZN(G1338GAT) );
  NOR2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U585 ( .A(G106GAT), .B(n521), .Z(n522) );
  XNOR2_X1 U586 ( .A(KEYINPUT44), .B(n522), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U588 ( .A(KEYINPUT110), .B(n525), .Z(n544) );
  NOR2_X1 U589 ( .A1(n544), .A2(n526), .ZN(n527) );
  XNOR2_X1 U590 ( .A(n527), .B(KEYINPUT111), .ZN(n528) );
  NOR2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n540) );
  NAND2_X1 U592 ( .A1(n540), .A2(n558), .ZN(n530) );
  XNOR2_X1 U593 ( .A(n530), .B(KEYINPUT112), .ZN(n531) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n531), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT49), .B(KEYINPUT114), .Z(n534) );
  INV_X1 U596 ( .A(n532), .ZN(n560) );
  NAND2_X1 U597 ( .A1(n540), .A2(n560), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(n536) );
  XOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT113), .Z(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n538) );
  NAND2_X1 U602 ( .A1(n540), .A2(n564), .ZN(n537) );
  XNOR2_X1 U603 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(G134GAT), .B(KEYINPUT51), .Z(n542) );
  NAND2_X1 U606 ( .A1(n540), .A2(n555), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(G1343GAT) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(KEYINPUT116), .ZN(n546) );
  INV_X1 U609 ( .A(n569), .ZN(n543) );
  NOR2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n554) );
  NAND2_X1 U611 ( .A1(n558), .A2(n554), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(G1344GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n548) );
  NAND2_X1 U614 ( .A1(n554), .A2(n560), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n548), .B(n547), .ZN(n550) );
  XOR2_X1 U616 ( .A(G148GAT), .B(KEYINPUT53), .Z(n549) );
  XNOR2_X1 U617 ( .A(n550), .B(n549), .ZN(G1345GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n552) );
  NAND2_X1 U619 ( .A1(n554), .A2(n579), .ZN(n551) );
  XNOR2_X1 U620 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n553), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT120), .ZN(n557) );
  XNOR2_X1 U624 ( .A(G162GAT), .B(n557), .ZN(G1347GAT) );
  NAND2_X1 U625 ( .A1(n565), .A2(n558), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n562) );
  NAND2_X1 U628 ( .A1(n565), .A2(n560), .ZN(n561) );
  XNOR2_X1 U629 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G176GAT), .ZN(G1349GAT) );
  NAND2_X1 U631 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n573) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n578) );
  NOR2_X1 U637 ( .A1(n571), .A2(n578), .ZN(n572) );
  XOR2_X1 U638 ( .A(n573), .B(n572), .Z(G1352GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n578), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT61), .B(KEYINPUT125), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(G204GAT), .B(n577), .Z(G1353GAT) );
  INV_X1 U643 ( .A(n578), .ZN(n583) );
  AND2_X1 U644 ( .A1(n579), .A2(n583), .ZN(n580) );
  XOR2_X1 U645 ( .A(KEYINPUT126), .B(n580), .Z(n581) );
  XNOR2_X1 U646 ( .A(G211GAT), .B(n581), .ZN(G1354GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n585) );
  NAND2_X1 U648 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

