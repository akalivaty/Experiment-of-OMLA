//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n562, new_n563, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1146, new_n1147, new_n1148;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  XNOR2_X1  g036(.A(KEYINPUT66), .B(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2105), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n467), .A2(G101), .A3(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT68), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n470), .A2(new_n467), .A3(G101), .A4(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT67), .B1(new_n473), .B2(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(KEYINPUT67), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(new_n476), .A3(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n473), .A2(KEYINPUT3), .ZN(new_n478));
  NAND3_X1  g053(.A1(new_n474), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n467), .A2(KEYINPUT66), .ZN(new_n480));
  INV_X1    g055(.A(KEYINPUT66), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G2105), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n480), .A2(new_n482), .A3(G137), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n472), .B1(new_n479), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT69), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n472), .B(new_n486), .C1(new_n479), .C2(new_n483), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n466), .B1(new_n485), .B2(new_n487), .ZN(G160));
  XNOR2_X1  g063(.A(new_n479), .B(KEYINPUT70), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(new_n467), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(G136), .ZN(new_n492));
  INV_X1    g067(.A(new_n462), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G124), .ZN(new_n496));
  OAI221_X1 g071(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n462), .C2(G112), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n492), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G162));
  NAND3_X1  g074(.A1(new_n480), .A2(new_n482), .A3(G138), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT4), .B1(new_n479), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n463), .A2(new_n462), .A3(new_n502), .A4(G138), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AND3_X1   g079(.A1(new_n474), .A2(new_n477), .A3(new_n478), .ZN(new_n505));
  AND2_X1   g080(.A1(G126), .A2(G2105), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n467), .A2(G114), .ZN(new_n507));
  OAI21_X1  g082(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n504), .A2(new_n510), .ZN(G164));
  XOR2_X1   g086(.A(KEYINPUT5), .B(G543), .Z(new_n512));
  AND2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g090(.A(KEYINPUT71), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n513), .A2(new_n514), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  XNOR2_X1  g093(.A(KEYINPUT5), .B(G543), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n517), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G88), .ZN(new_n523));
  NAND2_X1  g098(.A1(G75), .A2(G543), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT72), .ZN(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n512), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n515), .A2(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n527), .A2(G651), .B1(new_n529), .B2(G50), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n523), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  INV_X1    g107(.A(KEYINPUT74), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT7), .ZN(new_n535));
  INV_X1    g110(.A(G89), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n533), .B(new_n535), .C1(new_n521), .C2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n519), .A2(G63), .A3(G651), .ZN(new_n538));
  INV_X1    g113(.A(new_n529), .ZN(new_n539));
  XNOR2_X1  g114(.A(KEYINPUT73), .B(G51), .ZN(new_n540));
  OAI211_X1 g115(.A(new_n537), .B(new_n538), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n522), .A2(G89), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n533), .B1(new_n542), .B2(new_n535), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(G168));
  AOI22_X1  g119(.A1(new_n519), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n545));
  INV_X1    g120(.A(G651), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G52), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n547), .B1(new_n548), .B2(new_n539), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(new_n522), .B2(G90), .ZN(G171));
  XNOR2_X1  g125(.A(KEYINPUT76), .B(G81), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n522), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n519), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n553), .A2(new_n546), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n554), .A2(new_n555), .B1(G43), .B2(new_n529), .ZN(new_n556));
  OAI21_X1  g131(.A(KEYINPUT75), .B1(new_n553), .B2(new_n546), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n552), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  NAND4_X1  g135(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT8), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  NAND2_X1  g139(.A1(new_n529), .A2(G53), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT9), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n522), .A2(G91), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n519), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n566), .B(new_n567), .C1(new_n546), .C2(new_n568), .ZN(G299));
  INV_X1    g144(.A(G171), .ZN(G301));
  OR2_X1    g145(.A1(new_n541), .A2(new_n543), .ZN(G286));
  OR2_X1    g146(.A1(new_n519), .A2(G74), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G651), .B1(new_n529), .B2(G49), .ZN(new_n573));
  INV_X1    g148(.A(G87), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n521), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT77), .ZN(G288));
  AOI22_X1  g151(.A1(new_n519), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n577));
  OR2_X1    g152(.A1(new_n577), .A2(new_n546), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n516), .A2(new_n520), .A3(G86), .ZN(new_n579));
  OAI211_X1 g154(.A(G48), .B(G543), .C1(new_n513), .C2(new_n514), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT78), .ZN(new_n581));
  XNOR2_X1  g156(.A(new_n580), .B(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n578), .A2(new_n579), .A3(new_n582), .ZN(G305));
  NAND2_X1  g158(.A1(new_n529), .A2(G47), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n519), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI221_X1 g161(.A(new_n584), .B1(new_n546), .B2(new_n585), .C1(new_n521), .C2(new_n586), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT79), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n522), .A2(KEYINPUT10), .A3(G92), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  INV_X1    g166(.A(G92), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n521), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n512), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(new_n529), .B2(G54), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n589), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n589), .B1(new_n599), .B2(G868), .ZN(G321));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  NAND2_X1  g177(.A1(G299), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G168), .B2(new_n602), .ZN(G297));
  XOR2_X1   g179(.A(G297), .B(KEYINPUT80), .Z(G280));
  INV_X1    g180(.A(G559), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n599), .B1(new_n606), .B2(G860), .ZN(G148));
  NAND2_X1  g182(.A1(new_n558), .A2(new_n602), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n599), .A2(new_n606), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n602), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n491), .A2(G135), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n495), .A2(G123), .ZN(new_n613));
  OAI221_X1 g188(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n462), .C2(G111), .ZN(new_n614));
  AND3_X1   g189(.A1(new_n612), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(G2096), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(G2096), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n467), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n617), .A2(new_n618), .A3(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(G2427), .B(G2438), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2430), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT15), .B(G2435), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n627), .A2(KEYINPUT14), .A3(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(G1341), .B(G1348), .Z(new_n630));
  XNOR2_X1  g205(.A(G2443), .B(G2446), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n629), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2451), .B(G2454), .Z(new_n634));
  XNOR2_X1  g209(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n633), .A2(new_n636), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n637), .A2(G14), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT82), .Z(new_n640));
  INV_X1    g215(.A(new_n640), .ZN(G401));
  XNOR2_X1  g216(.A(G2067), .B(G2678), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2072), .B(G2078), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2084), .B(G2090), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT18), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(KEYINPUT17), .ZN(new_n648));
  OR2_X1    g223(.A1(new_n642), .A2(new_n645), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n645), .B1(new_n642), .B2(new_n643), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n650), .B1(new_n648), .B2(new_n642), .ZN(new_n651));
  INV_X1    g226(.A(KEYINPUT83), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  OAI221_X1 g229(.A(new_n647), .B1(new_n648), .B2(new_n649), .C1(new_n653), .C2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT84), .ZN(new_n656));
  XOR2_X1   g231(.A(G2096), .B(G2100), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(G227));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  AND2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT20), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n660), .A2(new_n663), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n660), .B2(new_n666), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G1991), .B(G1996), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(G1981), .B(G1986), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT85), .ZN(new_n673));
  XOR2_X1   g248(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n671), .B(new_n675), .ZN(G229));
  INV_X1    g251(.A(G29), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n677), .A2(G25), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n495), .A2(G119), .ZN(new_n679));
  OAI221_X1 g254(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n462), .C2(G107), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n491), .A2(G131), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n678), .B1(new_n684), .B2(new_n677), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT35), .B(G1991), .Z(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  MUX2_X1   g262(.A(G24), .B(G290), .S(G16), .Z(new_n688));
  OR2_X1    g263(.A1(new_n688), .A2(G1986), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(G1986), .ZN(new_n690));
  AND4_X1   g265(.A1(KEYINPUT88), .A2(new_n687), .A3(new_n689), .A4(new_n690), .ZN(new_n691));
  MUX2_X1   g266(.A(G23), .B(new_n575), .S(G16), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT33), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1976), .ZN(new_n694));
  INV_X1    g269(.A(G16), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G22), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT87), .Z(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(G303), .B2(G16), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(G1971), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n695), .A2(G6), .ZN(new_n700));
  INV_X1    g275(.A(G305), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n700), .B1(new_n701), .B2(new_n695), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT86), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT32), .B(G1981), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  NAND4_X1  g281(.A1(new_n694), .A2(new_n699), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  OR2_X1    g282(.A1(new_n707), .A2(KEYINPUT34), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(KEYINPUT34), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n691), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(KEYINPUT36), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n677), .A2(G32), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT26), .Z(new_n715));
  NAND3_X1  g290(.A1(new_n467), .A2(G105), .A3(G2104), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n495), .B2(G129), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT91), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(new_n491), .B2(G141), .ZN(new_n720));
  INV_X1    g295(.A(G141), .ZN(new_n721));
  NOR3_X1   g296(.A1(new_n490), .A2(KEYINPUT91), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n718), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n713), .B1(new_n724), .B2(new_n677), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT27), .B(G1996), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT92), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n725), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n677), .A2(G35), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G162), .B2(new_n677), .ZN(new_n730));
  INV_X1    g305(.A(G2090), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT94), .B(KEYINPUT29), .Z(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n728), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n736), .B1(new_n735), .B2(new_n733), .ZN(new_n737));
  NAND2_X1  g312(.A1(G299), .A2(G16), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n695), .A2(G20), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(KEYINPUT23), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1956), .ZN(new_n742));
  NOR2_X1   g317(.A1(G4), .A2(G16), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n599), .B2(G16), .ZN(new_n744));
  AOI21_X1  g319(.A(new_n742), .B1(G1348), .B2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n677), .A2(G26), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT28), .Z(new_n747));
  OAI221_X1 g322(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n462), .C2(G116), .ZN(new_n748));
  INV_X1    g323(.A(G140), .ZN(new_n749));
  INV_X1    g324(.A(G128), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n748), .B1(new_n490), .B2(new_n749), .C1(new_n750), .C2(new_n494), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n747), .B1(new_n751), .B2(G29), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G2067), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n677), .A2(G33), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT25), .Z(new_n756));
  AOI22_X1  g331(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n756), .B1(new_n462), .B2(new_n757), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G139), .B2(new_n491), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n754), .B1(new_n759), .B2(new_n677), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(G2072), .Z(new_n761));
  NAND3_X1  g336(.A1(new_n745), .A2(new_n753), .A3(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT24), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n677), .B1(new_n763), .B2(G34), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(KEYINPUT89), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(KEYINPUT89), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n763), .A2(G34), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n765), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(KEYINPUT90), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G160), .B2(G29), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2084), .ZN(new_n771));
  NOR2_X1   g346(.A1(G164), .A2(new_n677), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G27), .B2(new_n677), .ZN(new_n773));
  INV_X1    g348(.A(G2078), .ZN(new_n774));
  OR2_X1    g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n695), .A2(G5), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G171), .B2(new_n695), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n775), .B(new_n776), .C1(G1961), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n695), .A2(G19), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n559), .B2(new_n695), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(G1341), .Z(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G1348), .B2(new_n744), .ZN(new_n783));
  NOR4_X1   g358(.A1(new_n762), .A2(new_n771), .A3(new_n779), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n695), .A2(G21), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G168), .B2(new_n695), .ZN(new_n786));
  AND2_X1   g361(.A1(new_n786), .A2(G1966), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n778), .A2(G1961), .ZN(new_n788));
  INV_X1    g363(.A(G28), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n789), .A2(KEYINPUT30), .ZN(new_n790));
  AOI21_X1  g365(.A(G29), .B1(new_n789), .B2(KEYINPUT30), .ZN(new_n791));
  OR2_X1    g366(.A1(KEYINPUT31), .A2(G11), .ZN(new_n792));
  NAND2_X1  g367(.A1(KEYINPUT31), .A2(G11), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n790), .A2(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI211_X1 g369(.A(new_n788), .B(new_n794), .C1(new_n616), .C2(new_n677), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n786), .A2(G1966), .ZN(new_n796));
  OR3_X1    g371(.A1(new_n787), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n797), .A2(KEYINPUT93), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(KEYINPUT93), .ZN(new_n799));
  AND4_X1   g374(.A1(new_n737), .A2(new_n784), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n710), .A2(new_n711), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n712), .A2(new_n800), .A3(new_n801), .ZN(G150));
  XNOR2_X1  g377(.A(G150), .B(KEYINPUT95), .ZN(G311));
  NAND2_X1  g378(.A1(new_n599), .A2(G559), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT96), .B(KEYINPUT38), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n529), .A2(G55), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n519), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT97), .B(G93), .ZN(new_n809));
  OAI221_X1 g384(.A(new_n807), .B1(new_n546), .B2(new_n808), .C1(new_n521), .C2(new_n809), .ZN(new_n810));
  OR2_X1    g385(.A1(new_n558), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n558), .A2(new_n810), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n806), .B(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(KEYINPUT39), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n815), .A2(new_n816), .A3(G860), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n810), .A2(G860), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT37), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n817), .A2(new_n819), .ZN(G145));
  INV_X1    g395(.A(KEYINPUT99), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n723), .B(new_n759), .ZN(new_n822));
  OAI221_X1 g397(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n462), .C2(G118), .ZN(new_n823));
  INV_X1    g398(.A(G130), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n494), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G142), .B2(new_n491), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n620), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n822), .A2(new_n827), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT98), .ZN(new_n831));
  AND3_X1   g406(.A1(new_n501), .A2(new_n831), .A3(new_n503), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n831), .B1(new_n501), .B2(new_n503), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n510), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n751), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n751), .A2(new_n834), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n837), .A2(new_n684), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n835), .A2(new_n683), .A3(new_n836), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n830), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n498), .B(G160), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(new_n615), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n828), .A2(new_n838), .A3(new_n839), .A4(new_n829), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G37), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g422(.A(new_n843), .B1(new_n841), .B2(new_n844), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n821), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n848), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n850), .A2(KEYINPUT99), .A3(new_n846), .A4(new_n845), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(KEYINPUT100), .B(KEYINPUT40), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n852), .B(new_n853), .Z(G395));
  NAND2_X1  g429(.A1(new_n810), .A2(new_n602), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n813), .B(KEYINPUT101), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(new_n609), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n599), .B(G299), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT41), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n858), .B(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n857), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(G290), .B(G305), .ZN(new_n864));
  XNOR2_X1  g439(.A(G303), .B(new_n575), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(G290), .B(new_n701), .ZN(new_n867));
  INV_X1    g442(.A(new_n865), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  AND3_X1   g444(.A1(new_n866), .A2(new_n869), .A3(KEYINPUT102), .ZN(new_n870));
  AOI21_X1  g445(.A(KEYINPUT102), .B1(new_n866), .B2(new_n869), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n872), .A2(KEYINPUT42), .ZN(new_n873));
  AOI21_X1  g448(.A(KEYINPUT42), .B1(new_n866), .B2(new_n869), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT103), .ZN(new_n876));
  OAI211_X1 g451(.A(new_n860), .B(new_n863), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n863), .A2(new_n860), .ZN(new_n878));
  OAI211_X1 g453(.A(KEYINPUT103), .B(new_n878), .C1(new_n873), .C2(new_n874), .ZN(new_n879));
  AOI22_X1  g454(.A1(new_n877), .A2(new_n879), .B1(new_n876), .B2(new_n875), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n855), .B1(new_n880), .B2(new_n602), .ZN(G295));
  OAI21_X1  g456(.A(new_n855), .B1(new_n880), .B2(new_n602), .ZN(G331));
  NAND2_X1  g457(.A1(G286), .A2(G301), .ZN(new_n883));
  NAND2_X1  g458(.A1(G168), .A2(G171), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n813), .ZN(new_n886));
  INV_X1    g461(.A(new_n813), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n887), .A2(new_n883), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(new_n859), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(KEYINPUT105), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT105), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n887), .A2(new_n883), .A3(new_n892), .A4(new_n884), .ZN(new_n893));
  INV_X1    g468(.A(KEYINPUT104), .ZN(new_n894));
  AND3_X1   g469(.A1(new_n885), .A2(new_n894), .A3(new_n813), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n894), .B1(new_n885), .B2(new_n813), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n891), .B(new_n893), .C1(new_n895), .C2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n890), .B1(new_n897), .B2(new_n862), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n870), .A2(new_n871), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n846), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n898), .A2(new_n899), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(KEYINPUT43), .ZN(new_n904));
  AOI21_X1  g479(.A(G37), .B1(new_n898), .B2(new_n899), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n862), .A2(new_n889), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n897), .B2(new_n859), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(new_n872), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n905), .A2(KEYINPUT43), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g484(.A(KEYINPUT44), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n908), .A2(new_n900), .A3(new_n911), .A4(new_n846), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT106), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT43), .B1(new_n901), .B2(new_n902), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT106), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n905), .A2(new_n915), .A3(new_n911), .A4(new_n908), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT44), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n910), .A2(new_n919), .ZN(G397));
  XOR2_X1   g495(.A(new_n723), .B(G1996), .Z(new_n921));
  XOR2_X1   g496(.A(new_n751), .B(G2067), .Z(new_n922));
  AND2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n684), .A2(new_n686), .ZN(new_n924));
  OR2_X1    g499(.A1(new_n684), .A2(new_n686), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n923), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(G1384), .ZN(new_n928));
  AOI21_X1  g503(.A(KEYINPUT45), .B1(new_n834), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n466), .ZN(new_n930));
  INV_X1    g505(.A(new_n483), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n505), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n486), .B1(new_n932), .B2(new_n472), .ZN(new_n933));
  INV_X1    g508(.A(new_n487), .ZN(new_n934));
  OAI211_X1 g509(.A(G40), .B(new_n930), .C1(new_n933), .C2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n929), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n927), .A2(new_n937), .ZN(new_n938));
  NOR3_X1   g513(.A1(new_n937), .A2(G290), .A3(G1986), .ZN(new_n939));
  XNOR2_X1  g514(.A(new_n939), .B(KEYINPUT48), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n751), .A2(G2067), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n924), .B(KEYINPUT125), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n941), .B1(new_n942), .B2(new_n923), .ZN(new_n943));
  OAI22_X1  g518(.A1(new_n938), .A2(new_n940), .B1(new_n937), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n937), .B1(new_n922), .B2(new_n724), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT46), .B1(new_n937), .B2(G1996), .ZN(new_n946));
  OR3_X1    g521(.A1(new_n937), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n945), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT47), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n944), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G8), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n504), .A2(KEYINPUT98), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n501), .A2(new_n503), .A3(new_n831), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI21_X1  g529(.A(G1384), .B1(new_n954), .B2(new_n510), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n951), .B1(new_n955), .B2(new_n936), .ZN(new_n956));
  NAND2_X1  g531(.A1(G305), .A2(G1981), .ZN(new_n957));
  INV_X1    g532(.A(G1981), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n578), .A2(new_n579), .A3(new_n582), .A4(new_n958), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n957), .A2(KEYINPUT49), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT49), .B1(new_n957), .B2(new_n959), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI211_X1 g537(.A(G1976), .B(G288), .C1(new_n962), .C2(new_n956), .ZN(new_n963));
  INV_X1    g538(.A(new_n959), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n956), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n955), .A2(new_n936), .ZN(new_n966));
  OAI211_X1 g541(.A(new_n573), .B(G1976), .C1(new_n574), .C2(new_n521), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n966), .A2(G8), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT109), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n956), .A2(new_n970), .A3(new_n967), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(KEYINPUT52), .A3(new_n971), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n966), .A2(G8), .A3(new_n967), .ZN(new_n973));
  XNOR2_X1  g548(.A(KEYINPUT110), .B(G1976), .ZN(new_n974));
  AOI21_X1  g549(.A(KEYINPUT52), .B1(G288), .B2(new_n974), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n973), .A2(new_n975), .B1(new_n962), .B2(new_n956), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n972), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n978));
  OAI211_X1 g553(.A(G303), .B(G8), .C1(new_n978), .C2(KEYINPUT55), .ZN(new_n979));
  NOR2_X1   g554(.A1(G166), .A2(new_n951), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT108), .B(KEYINPUT55), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n504), .A2(new_n510), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n983), .A2(new_n928), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT50), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n834), .A2(new_n928), .ZN(new_n986));
  XNOR2_X1  g561(.A(KEYINPUT107), .B(KEYINPUT50), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n936), .B(new_n985), .C1(new_n986), .C2(new_n988), .ZN(new_n989));
  NOR2_X1   g564(.A1(new_n989), .A2(G2090), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT45), .B1(new_n983), .B2(new_n928), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n991), .A2(new_n935), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n834), .A2(KEYINPUT45), .A3(new_n928), .ZN(new_n993));
  AOI21_X1  g568(.A(G1971), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OAI211_X1 g569(.A(G8), .B(new_n982), .C1(new_n990), .C2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n965), .B1(new_n977), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT113), .ZN(new_n997));
  AND3_X1   g572(.A1(new_n995), .A2(new_n972), .A3(new_n976), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n986), .A2(new_n988), .ZN(new_n999));
  INV_X1    g574(.A(new_n984), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT50), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n935), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n999), .A2(new_n1002), .A3(new_n731), .ZN(new_n1003));
  OAI21_X1  g578(.A(KEYINPUT111), .B1(new_n1003), .B2(new_n994), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n992), .A2(new_n993), .ZN(new_n1005));
  INV_X1    g580(.A(G1971), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT111), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n999), .A2(new_n1002), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1007), .B(new_n1008), .C1(G2090), .C2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1004), .A2(G8), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n982), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n998), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n989), .A2(G2084), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n929), .B2(new_n935), .ZN(new_n1017));
  OAI211_X1 g592(.A(KEYINPUT112), .B(new_n936), .C1(new_n955), .C2(KEYINPUT45), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1000), .A2(KEYINPUT45), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G1966), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1015), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  NOR3_X1   g597(.A1(new_n1022), .A2(new_n951), .A3(G286), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n997), .B1(new_n1014), .B2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n998), .A2(new_n1013), .A3(new_n1023), .A4(KEYINPUT113), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT63), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1025), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n990), .B2(new_n994), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1027), .B1(new_n1029), .B2(new_n1012), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n998), .A2(new_n1023), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n996), .B1(new_n1028), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(G2078), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT119), .ZN(new_n1036));
  INV_X1    g611(.A(G1961), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n989), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1035), .A2(new_n1036), .A3(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n992), .A2(new_n993), .A3(new_n774), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n1033), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT120), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1040), .A2(KEYINPUT120), .A3(new_n1033), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1039), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1036), .B1(new_n1035), .B2(new_n1038), .ZN(new_n1047));
  OAI21_X1  g622(.A(G171), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT121), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  OAI211_X1 g625(.A(KEYINPUT121), .B(G171), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT62), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G168), .A2(new_n951), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n1022), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(KEYINPUT51), .B1(new_n1054), .B2(KEYINPUT118), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1055), .B(new_n1058), .C1(new_n1022), .C2(new_n951), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  AOI211_X1 g635(.A(new_n951), .B(new_n1058), .C1(new_n1022), .C2(G168), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n1053), .B(new_n1057), .C1(new_n1060), .C2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1014), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1052), .A2(new_n1062), .A3(KEYINPUT124), .A4(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1057), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1065), .A2(KEYINPUT62), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1058), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1015), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(G8), .B(new_n1068), .C1(new_n1071), .C2(G286), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1056), .B1(new_n1072), .B2(new_n1059), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1014), .B1(new_n1073), .B2(new_n1053), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT124), .B1(new_n1074), .B2(new_n1052), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1032), .B1(new_n1067), .B2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1047), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1077), .A2(G301), .A3(new_n1045), .A4(new_n1039), .ZN(new_n1078));
  INV_X1    g653(.A(new_n929), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1079), .A2(new_n936), .A3(new_n1034), .A4(new_n993), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1045), .A2(new_n1038), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT122), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1081), .A2(new_n1082), .A3(G171), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1038), .A2(new_n1080), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT122), .B1(new_n1085), .B2(G301), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1078), .A2(new_n1083), .A3(new_n1086), .A4(KEYINPUT54), .ZN(new_n1087));
  AND3_X1   g662(.A1(new_n1087), .A2(new_n1065), .A3(new_n1063), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1085), .A2(G301), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1050), .A2(new_n1051), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1092), .A3(KEYINPUT123), .ZN(new_n1093));
  INV_X1    g668(.A(G1956), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1009), .A2(new_n1094), .ZN(new_n1095));
  XNOR2_X1  g670(.A(KEYINPUT56), .B(G2072), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n992), .A2(new_n993), .A3(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT114), .B(KEYINPUT57), .ZN(new_n1098));
  XNOR2_X1  g673(.A(G299), .B(new_n1098), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1095), .A2(new_n1097), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT115), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1099), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1102), .B2(new_n1101), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n966), .A2(G2067), .ZN(new_n1105));
  INV_X1    g680(.A(G1348), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(new_n989), .ZN(new_n1107));
  INV_X1    g682(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n599), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1100), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1107), .B(new_n599), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT60), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1101), .B(new_n1099), .ZN(new_n1113));
  OAI22_X1  g688(.A1(new_n1111), .A2(new_n1112), .B1(new_n1113), .B2(KEYINPUT61), .ZN(new_n1114));
  XOR2_X1   g689(.A(KEYINPUT58), .B(G1341), .Z(new_n1115));
  NAND2_X1  g690(.A1(new_n966), .A2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n1005), .B2(G1996), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1117), .A2(new_n559), .ZN(new_n1118));
  XNOR2_X1  g693(.A(KEYINPUT116), .B(KEYINPUT59), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1107), .A2(new_n1112), .A3(new_n599), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1114), .A2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(new_n1100), .B(KEYINPUT117), .Z(new_n1125));
  NAND3_X1  g700(.A1(new_n1125), .A2(KEYINPUT61), .A3(new_n1104), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1110), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1088), .A2(new_n1092), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT123), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1127), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1076), .B1(new_n1093), .B2(new_n1130), .ZN(new_n1131));
  XOR2_X1   g706(.A(G290), .B(G1986), .Z(new_n1132));
  AOI21_X1  g707(.A(new_n937), .B1(new_n927), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n950), .B1(new_n1131), .B2(new_n1133), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g709(.A1(G229), .A2(G227), .A3(new_n460), .ZN(new_n1136));
  NAND2_X1  g710(.A1(new_n1136), .A2(new_n640), .ZN(new_n1137));
  NAND2_X1  g711(.A1(new_n1137), .A2(KEYINPUT126), .ZN(new_n1138));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n1139));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n1139), .A3(new_n640), .ZN(new_n1140));
  AOI22_X1  g714(.A1(new_n849), .A2(new_n851), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g715(.A(KEYINPUT127), .ZN(new_n1142));
  AND3_X1   g716(.A1(new_n917), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g717(.A(new_n1142), .B1(new_n917), .B2(new_n1141), .ZN(new_n1144));
  NOR2_X1   g718(.A1(new_n1143), .A2(new_n1144), .ZN(G308));
  NAND2_X1  g719(.A1(new_n917), .A2(new_n1141), .ZN(new_n1146));
  NAND2_X1  g720(.A1(new_n1146), .A2(KEYINPUT127), .ZN(new_n1147));
  NAND3_X1  g721(.A1(new_n917), .A2(new_n1141), .A3(new_n1142), .ZN(new_n1148));
  NAND2_X1  g722(.A1(new_n1147), .A2(new_n1148), .ZN(G225));
endmodule


