//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 0 0 1 0 1 0 0 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 1 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 1 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  XOR2_X1   g003(.A(G119), .B(G128), .Z(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT24), .B(G110), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT23), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G128), .ZN(new_n195));
  INV_X1    g009(.A(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT23), .A3(G119), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n195), .B(new_n197), .C1(G119), .C2(new_n196), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G110), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT72), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(KEYINPUT72), .A3(G110), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n192), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT73), .B(G125), .ZN(new_n204));
  OR2_X1    g018(.A1(KEYINPUT16), .A2(G140), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OR2_X1    g020(.A1(G125), .A2(G140), .ZN(new_n207));
  INV_X1    g021(.A(G140), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n204), .B2(new_n208), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n206), .B1(new_n209), .B2(KEYINPUT16), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G146), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  AOI211_X1 g026(.A(new_n212), .B(new_n206), .C1(KEYINPUT16), .C2(new_n209), .ZN(new_n213));
  OAI21_X1  g027(.A(new_n203), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT74), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(G146), .ZN(new_n216));
  XNOR2_X1  g030(.A(G125), .B(G140), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n212), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n190), .A2(new_n191), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n219), .B1(new_n198), .B2(G110), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n216), .A2(new_n218), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n214), .A2(new_n215), .A3(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT22), .B(G137), .ZN(new_n223));
  INV_X1    g037(.A(G953), .ZN(new_n224));
  AND3_X1   g038(.A1(new_n224), .A2(G221), .A3(G234), .ZN(new_n225));
  XOR2_X1   g039(.A(new_n223), .B(new_n225), .Z(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n222), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n214), .A2(new_n221), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT74), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n222), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n228), .B1(new_n231), .B2(new_n226), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT25), .B1(new_n232), .B2(new_n188), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n214), .A2(new_n215), .A3(new_n221), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n215), .B1(new_n214), .B2(new_n221), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n226), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n222), .A2(new_n227), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n236), .A2(new_n188), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT25), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n189), .B1(new_n233), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n189), .A2(G902), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n232), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT32), .ZN(new_n245));
  XNOR2_X1  g059(.A(KEYINPUT2), .B(G113), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(G116), .B(G119), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n248), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n246), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n212), .A2(G143), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n253), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(G143), .B(G146), .ZN(new_n260));
  INV_X1    g074(.A(new_n258), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(KEYINPUT65), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n259), .A2(new_n262), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n255), .A2(KEYINPUT64), .A3(G146), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT64), .B1(new_n255), .B2(G146), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n254), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G137), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n270), .A2(G134), .B1(KEYINPUT66), .B2(KEYINPUT11), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(G134), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(G131), .ZN(new_n274));
  INV_X1    g088(.A(G134), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(G137), .ZN(new_n276));
  NAND2_X1  g090(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(KEYINPUT66), .A2(KEYINPUT11), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n276), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AND3_X1   g094(.A1(new_n273), .A2(new_n274), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n274), .B1(new_n273), .B2(new_n280), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n263), .B(new_n269), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT30), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT1), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n260), .A2(new_n285), .A3(G128), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT64), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n287), .B1(new_n212), .B2(G143), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n255), .A2(KEYINPUT64), .A3(G146), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n288), .A2(new_n289), .B1(G143), .B2(new_n212), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n285), .B1(G143), .B2(new_n212), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n291), .A2(new_n196), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n286), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n273), .A2(new_n274), .A3(new_n280), .ZN(new_n294));
  OAI21_X1  g108(.A(G131), .B1(new_n276), .B2(new_n272), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n293), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n283), .A2(new_n284), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n284), .B1(new_n283), .B2(new_n296), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n252), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n252), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n283), .A2(new_n300), .A3(new_n296), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT26), .B(G101), .ZN(new_n302));
  NOR2_X1   g116(.A1(G237), .A2(G953), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G210), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n302), .B(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT67), .B(KEYINPUT27), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n305), .A2(new_n306), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n299), .A2(new_n301), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT31), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n299), .A2(KEYINPUT31), .A3(new_n301), .A4(new_n310), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n301), .A2(KEYINPUT69), .A3(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(KEYINPUT69), .B1(new_n301), .B2(new_n315), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n283), .A2(new_n300), .A3(new_n296), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n300), .B1(new_n283), .B2(new_n296), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT28), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n319), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT68), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n308), .B2(new_n309), .ZN(new_n325));
  INV_X1    g139(.A(new_n309), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT68), .A3(new_n307), .ZN(new_n327));
  AND2_X1   g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n313), .A2(new_n314), .B1(new_n323), .B2(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(G472), .A2(G902), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n245), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n313), .A2(new_n314), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n323), .A2(new_n329), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n336), .A2(KEYINPUT32), .A3(new_n331), .ZN(new_n337));
  AND2_X1   g151(.A1(new_n333), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT69), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n339), .B1(new_n320), .B2(KEYINPUT28), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n322), .A2(new_n340), .A3(new_n316), .A4(new_n328), .ZN(new_n341));
  INV_X1    g155(.A(new_n310), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n281), .A2(new_n282), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n263), .A2(new_n269), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n296), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT30), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n283), .A2(new_n284), .A3(new_n296), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n300), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n342), .B1(new_n348), .B2(new_n320), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT29), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n341), .A2(new_n349), .A3(KEYINPUT70), .A4(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n342), .A2(new_n350), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n294), .A2(new_n295), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n270), .A2(G134), .ZN(new_n354));
  INV_X1    g168(.A(new_n279), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n354), .B1(new_n355), .B2(new_n277), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n275), .A2(G137), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n357), .B1(new_n276), .B2(new_n278), .ZN(new_n358));
  OAI21_X1  g172(.A(G131), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n294), .ZN(new_n360));
  AOI22_X1  g174(.A1(new_n259), .A2(new_n262), .B1(new_n266), .B2(new_n268), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n293), .A2(new_n353), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT71), .B1(new_n362), .B2(new_n300), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n345), .A2(new_n252), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n301), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n363), .B1(new_n365), .B2(KEYINPUT71), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n319), .B(new_n352), .C1(new_n366), .C2(new_n315), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n351), .A2(new_n188), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n299), .A2(new_n301), .ZN(new_n369));
  AOI21_X1  g183(.A(KEYINPUT29), .B1(new_n369), .B2(new_n342), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT70), .B1(new_n370), .B2(new_n341), .ZN(new_n371));
  OAI21_X1  g185(.A(G472), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n244), .B1(new_n338), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT75), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n375));
  INV_X1    g189(.A(new_n292), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n266), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n375), .B1(new_n377), .B2(new_n286), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n379), .A2(G104), .ZN(new_n380));
  INV_X1    g194(.A(G104), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n381), .A2(G107), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT76), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n383), .A2(KEYINPUT3), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n380), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n379), .A2(G104), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT3), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(KEYINPUT76), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n383), .A2(KEYINPUT3), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n386), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(G101), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT78), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n381), .A2(G107), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n391), .B1(new_n394), .B2(new_n386), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n392), .A2(new_n393), .A3(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n393), .B1(new_n392), .B2(new_n396), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n378), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n286), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n196), .B1(new_n291), .B2(KEYINPUT77), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n254), .A2(KEYINPUT1), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT77), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n400), .B1(new_n405), .B2(new_n257), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n392), .A2(new_n396), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n375), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n391), .B1(new_n385), .B2(new_n390), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT4), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n392), .A2(KEYINPUT4), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n411), .B(new_n361), .C1(new_n412), .C2(new_n409), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT79), .B1(new_n281), .B2(new_n282), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT79), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n359), .A2(new_n415), .A3(new_n294), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n399), .A2(new_n408), .A3(new_n413), .A4(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT81), .ZN(new_n419));
  XNOR2_X1  g233(.A(G110), .B(G140), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n224), .A2(G227), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n420), .B(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n418), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n399), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n408), .A2(new_n413), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n360), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n419), .B1(new_n418), .B2(new_n423), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT12), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n406), .A2(new_n407), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n387), .A2(KEYINPUT76), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n382), .B1(new_n384), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n394), .B1(new_n388), .B2(new_n386), .ZN(new_n435));
  NOR3_X1   g249(.A1(new_n434), .A2(new_n435), .A3(G101), .ZN(new_n436));
  OAI21_X1  g250(.A(KEYINPUT78), .B1(new_n436), .B2(new_n395), .ZN(new_n437));
  INV_X1    g251(.A(new_n293), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n392), .A2(new_n393), .A3(new_n396), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n432), .B1(new_n440), .B2(KEYINPUT80), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT80), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n437), .A2(new_n442), .A3(new_n438), .A4(new_n439), .ZN(new_n443));
  AOI211_X1 g257(.A(new_n431), .B(new_n343), .C1(new_n441), .C2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(KEYINPUT80), .ZN(new_n445));
  INV_X1    g259(.A(new_n432), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT12), .B1(new_n447), .B2(new_n360), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n418), .B1(new_n444), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n430), .B1(new_n449), .B2(new_n422), .ZN(new_n450));
  OAI21_X1  g264(.A(G469), .B1(new_n450), .B2(G902), .ZN(new_n451));
  XOR2_X1   g265(.A(KEYINPUT82), .B(G469), .Z(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n418), .A2(new_n423), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n447), .A2(new_n360), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n431), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n447), .A2(KEYINPUT12), .A3(new_n360), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n454), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n423), .B1(new_n427), .B2(new_n418), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n188), .B(new_n453), .C1(new_n458), .C2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n451), .A2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT9), .B(G234), .ZN(new_n462));
  OAI21_X1  g276(.A(G221), .B1(new_n462), .B2(G902), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n303), .A2(G143), .A3(G214), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(G143), .B1(new_n303), .B2(G214), .ZN(new_n467));
  OAI21_X1  g281(.A(G131), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(G237), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n224), .A3(G214), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(new_n255), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(new_n274), .A3(new_n465), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT19), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n217), .A2(new_n474), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n212), .B(new_n475), .C1(new_n209), .C2(new_n474), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n216), .A2(new_n473), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(G113), .B(G122), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n478), .B(G104), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g294(.A(KEYINPUT91), .B(new_n218), .C1(new_n209), .C2(new_n212), .ZN(new_n481));
  NAND2_X1  g295(.A1(KEYINPUT18), .A2(G131), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n482), .B1(new_n466), .B2(new_n467), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n471), .A2(KEYINPUT18), .A3(G131), .A4(new_n465), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(KEYINPUT73), .B(G125), .Z(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(G140), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT91), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n487), .A2(new_n488), .A3(G146), .A4(new_n207), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n481), .A2(new_n485), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(KEYINPUT92), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n481), .A2(new_n485), .A3(new_n489), .A4(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n480), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(G475), .A2(G902), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n211), .A2(new_n213), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT17), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n468), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n468), .A2(new_n498), .A3(new_n472), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n497), .A2(new_n501), .B1(new_n491), .B2(new_n493), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n495), .B(new_n496), .C1(new_n502), .C2(new_n479), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT20), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n497), .A2(new_n501), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(new_n494), .ZN(new_n506));
  INV_X1    g320(.A(new_n479), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT20), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n508), .A2(new_n509), .A3(new_n495), .A4(new_n496), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n507), .A2(KEYINPUT93), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n506), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n502), .A2(new_n512), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(new_n188), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G475), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT94), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n504), .A2(new_n510), .B1(new_n516), .B2(G475), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT94), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G952), .ZN(new_n524));
  AOI211_X1 g338(.A(G953), .B(new_n524), .C1(G234), .C2(G237), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n188), .B(new_n224), .C1(G234), .C2(G237), .ZN(new_n526));
  XNOR2_X1  g340(.A(KEYINPUT21), .B(G898), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT95), .B(G122), .ZN(new_n530));
  INV_X1    g344(.A(G116), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(G122), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n532), .B(new_n379), .C1(G116), .C2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(G128), .B(G143), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n535), .B(new_n275), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT14), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n533), .A2(G116), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n532), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n538), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT96), .ZN(new_n542));
  OAI21_X1  g356(.A(G107), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n537), .A2(new_n543), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n462), .A2(new_n187), .A3(G953), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT97), .ZN(new_n546));
  NOR2_X1   g360(.A1(new_n530), .A2(new_n531), .ZN(new_n547));
  OAI21_X1  g361(.A(G107), .B1(new_n547), .B2(new_n539), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n534), .A2(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT13), .B1(new_n196), .B2(G143), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(new_n275), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n551), .B(new_n535), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  AND3_X1   g367(.A1(new_n544), .A2(new_n546), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n546), .B1(new_n544), .B2(new_n553), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n188), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G478), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n557), .A2(KEYINPUT15), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI221_X1 g373(.A(new_n188), .B1(KEYINPUT15), .B2(new_n557), .C1(new_n554), .C2(new_n555), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n523), .A2(new_n529), .A3(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n464), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n411), .B(new_n252), .C1(new_n412), .C2(new_n409), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT83), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n437), .A2(new_n439), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT5), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(new_n194), .A3(G116), .ZN(new_n569));
  OAI211_X1 g383(.A(G113), .B(new_n569), .C1(new_n250), .C2(new_n568), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n570), .A2(new_n249), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n566), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n249), .ZN(new_n573));
  AOI211_X1 g387(.A(KEYINPUT83), .B(new_n573), .C1(new_n437), .C2(new_n439), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n565), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(G110), .B(G122), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n576), .B(new_n565), .C1(new_n572), .C2(new_n574), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(KEYINPUT6), .A3(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n377), .A2(KEYINPUT84), .A3(new_n286), .A4(new_n204), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n204), .B1(new_n263), .B2(new_n269), .ZN(new_n582));
  OAI211_X1 g396(.A(new_n286), .B(new_n204), .C1(new_n290), .C2(new_n292), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT84), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n581), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT85), .B(G224), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n587), .A2(G953), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n586), .B(new_n588), .Z(new_n589));
  INV_X1    g403(.A(KEYINPUT6), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n575), .A2(new_n590), .A3(new_n577), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n580), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(KEYINPUT86), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT86), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n580), .A2(new_n594), .A3(new_n589), .A4(new_n591), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT7), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n588), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  AND2_X1   g413(.A1(KEYINPUT88), .A2(KEYINPUT7), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  AND3_X1   g415(.A1(new_n586), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n599), .B1(new_n586), .B2(new_n601), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n570), .A2(KEYINPUT87), .A3(new_n249), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT87), .B1(new_n570), .B2(new_n249), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n606), .A2(new_n567), .B1(new_n573), .B2(new_n407), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n576), .B(KEYINPUT8), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  OAI22_X1  g423(.A1(new_n602), .A2(new_n603), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT89), .ZN(new_n611));
  OAI21_X1  g425(.A(new_n579), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n603), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n586), .A2(new_n599), .A3(new_n601), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  OR2_X1    g429(.A1(new_n604), .A2(new_n605), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n397), .A2(new_n398), .ZN(new_n617));
  INV_X1    g431(.A(new_n407), .ZN(new_n618));
  OAI22_X1  g432(.A1(new_n616), .A2(new_n617), .B1(new_n571), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(new_n608), .ZN(new_n620));
  AOI21_X1  g434(.A(KEYINPUT89), .B1(new_n615), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n188), .B1(new_n612), .B2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n596), .A2(new_n623), .ZN(new_n624));
  OAI21_X1  g438(.A(G210), .B1(G237), .B2(G902), .ZN(new_n625));
  INV_X1    g439(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n624), .A2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT90), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n596), .A2(new_n625), .A3(new_n623), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(G214), .B1(G237), .B2(G902), .ZN(new_n631));
  AOI211_X1 g445(.A(new_n626), .B(new_n622), .C1(new_n593), .C2(new_n595), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(KEYINPUT90), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n564), .A2(new_n630), .A3(new_n631), .A4(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n374), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n391), .ZN(G3));
  AOI21_X1  g450(.A(new_n625), .B1(new_n596), .B2(new_n623), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n631), .B1(new_n637), .B2(new_n632), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n640));
  INV_X1    g454(.A(G472), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n336), .B(new_n188), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  OAI211_X1 g456(.A(KEYINPUT98), .B(G472), .C1(new_n330), .C2(G902), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n642), .A2(new_n643), .A3(new_n241), .A4(new_n243), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n464), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n511), .A2(new_n521), .A3(new_n517), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n521), .B1(new_n511), .B2(new_n517), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT33), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n649), .B1(new_n554), .B2(new_n555), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT99), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n554), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n555), .A2(KEYINPUT100), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT100), .ZN(new_n655));
  AOI22_X1  g469(.A1(new_n537), .A2(new_n543), .B1(new_n549), .B2(new_n552), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n655), .B1(new_n656), .B2(new_n546), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n653), .A2(new_n654), .A3(KEYINPUT33), .A4(new_n657), .ZN(new_n658));
  OAI211_X1 g472(.A(KEYINPUT99), .B(new_n649), .C1(new_n554), .C2(new_n555), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n557), .A2(G902), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n652), .A2(new_n658), .A3(new_n659), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n556), .A2(new_n557), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n648), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n664), .A2(new_n528), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n639), .A2(new_n645), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT34), .B(G104), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G6));
  NAND4_X1  g482(.A1(new_n511), .A2(new_n561), .A3(new_n529), .A4(new_n517), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(new_n671));
  OAI211_X1 g485(.A(new_n671), .B(new_n631), .C1(new_n637), .C2(new_n632), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n645), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT35), .B(G107), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  AND2_X1   g490(.A1(new_n642), .A2(new_n643), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n227), .A2(KEYINPUT36), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n229), .B(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n242), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n241), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n634), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT37), .B(G110), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  NAND3_X1  g499(.A1(new_n372), .A2(new_n337), .A3(new_n333), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n686), .A2(new_n461), .A3(new_n463), .A4(new_n681), .ZN(new_n687));
  INV_X1    g501(.A(G900), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n526), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n525), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n520), .A2(new_n561), .A3(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n638), .A2(new_n687), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n196), .ZN(G30));
  NAND2_X1  g508(.A1(new_n630), .A2(new_n633), .ZN(new_n695));
  XNOR2_X1  g509(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n696));
  INV_X1    g510(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n630), .A2(new_n633), .A3(new_n696), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n523), .A2(new_n562), .ZN(new_n700));
  INV_X1    g514(.A(new_n681), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n311), .B1(new_n366), .B2(new_n328), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n702), .A2(new_n188), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n333), .B(new_n337), .C1(new_n641), .C2(new_n703), .ZN(new_n704));
  AND4_X1   g518(.A1(new_n631), .A2(new_n700), .A3(new_n701), .A4(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n698), .A2(new_n699), .A3(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT103), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n698), .A2(new_n708), .A3(new_n699), .A4(new_n705), .ZN(new_n709));
  INV_X1    g523(.A(new_n464), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n691), .B(KEYINPUT39), .ZN(new_n711));
  AND2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT40), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n707), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G143), .ZN(G45));
  NOR2_X1   g529(.A1(new_n638), .A2(new_n687), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n519), .A2(new_n522), .A3(new_n663), .A4(new_n691), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G146), .ZN(G48));
  INV_X1    g534(.A(G469), .ZN(new_n721));
  INV_X1    g535(.A(new_n454), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n722), .B1(new_n444), .B2(new_n448), .ZN(new_n723));
  INV_X1    g537(.A(new_n459), .ZN(new_n724));
  AOI21_X1  g538(.A(G902), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI211_X1 g539(.A(new_n460), .B(new_n463), .C1(new_n721), .C2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT104), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n723), .A2(new_n724), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n188), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(G469), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n731), .A2(KEYINPUT104), .A3(new_n463), .A4(new_n460), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n189), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n232), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n238), .A2(new_n239), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n737), .B1(new_n232), .B2(new_n242), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n686), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n733), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n740), .A2(new_n639), .A3(new_n665), .ZN(new_n741));
  XNOR2_X1  g555(.A(KEYINPUT41), .B(G113), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(KEYINPUT105), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n741), .B(new_n743), .ZN(G15));
  AOI21_X1  g558(.A(KEYINPUT106), .B1(new_n673), .B2(new_n740), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  NOR4_X1   g560(.A1(new_n672), .A2(new_n733), .A3(new_n746), .A4(new_n739), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n531), .ZN(G18));
  NOR2_X1   g563(.A1(new_n638), .A2(new_n733), .ZN(new_n750));
  INV_X1    g564(.A(new_n563), .ZN(new_n751));
  AND2_X1   g565(.A1(new_n686), .A2(new_n681), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n750), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G119), .ZN(G21));
  NOR2_X1   g568(.A1(new_n733), .A2(new_n528), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT71), .B1(new_n320), .B2(new_n321), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT71), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n301), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n315), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n340), .A2(new_n316), .ZN(new_n760));
  OAI21_X1  g574(.A(KEYINPUT107), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT107), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n762), .B(new_n319), .C1(new_n366), .C2(new_n315), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n761), .A2(new_n763), .A3(new_n329), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n334), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(new_n331), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n336), .A2(new_n188), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n766), .A2(KEYINPUT108), .B1(G472), .B2(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n765), .A2(new_n769), .A3(new_n331), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(new_n738), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n755), .A2(new_n639), .A3(new_n772), .A4(new_n700), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G122), .ZN(G24));
  AND2_X1   g588(.A1(new_n313), .A2(new_n314), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n319), .B1(new_n366), .B2(new_n315), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n328), .B1(new_n776), .B2(KEYINPUT107), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n775), .B1(new_n777), .B2(new_n763), .ZN(new_n778));
  OAI21_X1  g592(.A(KEYINPUT108), .B1(new_n778), .B2(new_n332), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n767), .A2(G472), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n779), .A2(new_n681), .A3(new_n770), .A4(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT109), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n768), .A2(KEYINPUT109), .A3(new_n681), .A4(new_n770), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n648), .A2(KEYINPUT110), .A3(new_n663), .A4(new_n691), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT110), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n717), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n785), .A2(new_n750), .A3(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G125), .ZN(G27));
  INV_X1    g606(.A(new_n631), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n793), .B1(new_n630), .B2(new_n633), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n794), .A2(new_n373), .A3(new_n710), .A4(new_n790), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT42), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI211_X1 g611(.A(new_n793), .B(new_n464), .C1(new_n630), .C2(new_n633), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(KEYINPUT42), .A3(new_n373), .A4(new_n790), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G131), .ZN(G33));
  INV_X1    g615(.A(new_n692), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n794), .A2(new_n373), .A3(new_n710), .A4(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G134), .ZN(G36));
  NOR2_X1   g618(.A1(new_n677), .A2(new_n701), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n523), .A2(new_n663), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT43), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT43), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n523), .A2(new_n808), .A3(new_n663), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n805), .A2(new_n807), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT112), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT44), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n811), .B1(new_n810), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n810), .A2(new_n812), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n695), .A2(new_n631), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT111), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n463), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n450), .A2(KEYINPUT45), .ZN(new_n820));
  OAI21_X1  g634(.A(G469), .B1(new_n450), .B2(KEYINPUT45), .ZN(new_n821));
  OAI22_X1  g635(.A1(new_n820), .A2(new_n821), .B1(new_n721), .B2(new_n188), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT46), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n822), .A2(new_n823), .B1(new_n725), .B2(new_n453), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n819), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n826), .A2(new_n711), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n794), .B(new_n828), .C1(new_n812), .C2(new_n810), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n815), .A2(new_n818), .A3(new_n827), .A4(new_n829), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n830), .B(G137), .ZN(G39));
  NOR3_X1   g645(.A1(new_n738), .A2(new_n686), .A3(new_n717), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n826), .A2(KEYINPUT47), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n826), .A2(KEYINPUT47), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n794), .B(new_n832), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G140), .ZN(G42));
  AOI21_X1  g651(.A(new_n789), .B1(new_n783), .B2(new_n784), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n710), .A3(new_n794), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n520), .A2(new_n562), .A3(new_n691), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n794), .A2(new_n710), .A3(new_n752), .A4(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n803), .A2(new_n839), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n634), .B1(new_n374), .B2(new_n682), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n748), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n519), .A2(new_n522), .A3(new_n662), .A4(new_n661), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n562), .B1(new_n646), .B2(new_n647), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n845), .A2(new_n846), .A3(new_n529), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n847), .A2(new_n464), .A3(new_n644), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(new_n631), .A3(new_n633), .A4(new_n630), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n741), .A2(new_n849), .A3(new_n773), .A4(new_n753), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n800), .A2(new_n842), .A3(new_n844), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n716), .A2(new_n802), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n701), .A2(new_n691), .A3(new_n704), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n639), .A2(new_n710), .A3(new_n700), .A4(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n791), .A2(new_n852), .A3(new_n719), .A4(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(KEYINPUT52), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n693), .B1(new_n838), .B2(new_n750), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n858), .A3(new_n719), .A4(new_n854), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT116), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n856), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n851), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT53), .ZN(new_n865));
  AND4_X1   g679(.A1(new_n800), .A2(new_n842), .A3(new_n844), .A4(new_n850), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n791), .A2(new_n852), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT52), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n856), .A2(new_n859), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n866), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n865), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT54), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n866), .A2(KEYINPUT53), .A3(new_n869), .ZN(new_n876));
  OAI211_X1 g690(.A(new_n875), .B(new_n876), .C1(new_n864), .C2(KEYINPUT53), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n807), .A2(new_n525), .A3(new_n809), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n771), .ZN(new_n880));
  OR3_X1    g694(.A1(new_n733), .A2(KEYINPUT119), .A3(new_n631), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT119), .B1(new_n733), .B2(new_n631), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n880), .A2(new_n881), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n698), .A2(new_n699), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT50), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT50), .B1(new_n883), .B2(new_n884), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n704), .A2(new_n244), .A3(new_n690), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n794), .A2(new_n728), .A3(new_n732), .A4(new_n890), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n891), .A2(new_n648), .A3(new_n663), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n817), .A2(new_n733), .A3(new_n879), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n892), .B1(new_n785), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT51), .ZN(new_n895));
  INV_X1    g709(.A(new_n835), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n731), .A2(new_n460), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n819), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n896), .A2(new_n833), .A3(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n880), .A2(new_n794), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n895), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n889), .A2(new_n894), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT120), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT120), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n889), .A2(new_n901), .A3(new_n904), .A4(new_n894), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n896), .A2(new_n833), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n898), .B(KEYINPUT117), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n900), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(KEYINPUT118), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n889), .A2(new_n910), .A3(new_n894), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n909), .A2(KEYINPUT118), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n895), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n893), .A2(new_n373), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT48), .Z(new_n915));
  AOI211_X1 g729(.A(new_n524), .B(G953), .C1(new_n880), .C2(new_n750), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(new_n891), .B2(new_n664), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n906), .A2(new_n913), .A3(new_n918), .ZN(new_n919));
  OAI22_X1  g733(.A1(new_n878), .A2(new_n919), .B1(G952), .B2(G953), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT49), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n897), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n738), .A2(new_n631), .A3(new_n463), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n923), .A2(KEYINPUT113), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(KEYINPUT113), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n806), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n922), .B1(new_n927), .B2(KEYINPUT114), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(KEYINPUT114), .B2(new_n927), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n929), .B(KEYINPUT115), .Z(new_n930));
  AOI21_X1  g744(.A(new_n704), .B1(new_n897), .B2(new_n921), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n884), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n920), .A2(new_n932), .ZN(G75));
  OAI21_X1  g747(.A(new_n876), .B1(new_n864), .B2(KEYINPUT53), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n934), .A2(G210), .A3(G902), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT56), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n580), .A2(new_n591), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n589), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT55), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n935), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n939), .B1(new_n935), .B2(new_n936), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n224), .A2(G952), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(G51));
  NOR2_X1   g757(.A1(new_n721), .A2(new_n188), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n944), .B(KEYINPUT57), .ZN(new_n945));
  AND3_X1   g759(.A1(new_n856), .A2(new_n859), .A3(new_n862), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n862), .B1(new_n856), .B2(new_n859), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n871), .B1(new_n948), .B2(new_n851), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n875), .B1(new_n949), .B2(new_n876), .ZN(new_n950));
  INV_X1    g764(.A(new_n877), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n945), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n729), .B(KEYINPUT121), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n934), .A2(G902), .ZN(new_n955));
  OR3_X1    g769(.A1(new_n955), .A2(new_n820), .A3(new_n821), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n942), .B1(new_n954), .B2(new_n956), .ZN(G54));
  NAND2_X1  g771(.A1(KEYINPUT58), .A2(G475), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n508), .ZN(new_n960));
  INV_X1    g774(.A(new_n495), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n959), .A2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n942), .ZN(new_n964));
  OAI22_X1  g778(.A1(new_n955), .A2(new_n958), .B1(new_n960), .B2(new_n961), .ZN(new_n965));
  AND3_X1   g779(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(G60));
  NAND3_X1  g780(.A1(new_n652), .A2(new_n658), .A3(new_n659), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(G478), .A2(G902), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT59), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n968), .B1(new_n878), .B2(new_n970), .ZN(new_n971));
  AND2_X1   g785(.A1(new_n968), .A2(new_n970), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(new_n950), .B2(new_n951), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n964), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n971), .A2(new_n974), .ZN(G63));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(KEYINPUT60), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n934), .A2(new_n679), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n964), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n232), .B1(new_n934), .B2(new_n979), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n976), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT122), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n978), .B1(new_n949), .B2(new_n876), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(new_n232), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n982), .A2(KEYINPUT122), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n980), .A2(KEYINPUT61), .A3(new_n964), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n983), .B1(new_n988), .B2(new_n989), .ZN(G66));
  OAI21_X1  g804(.A(G953), .B1(new_n587), .B2(new_n527), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n844), .A2(new_n850), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n991), .B1(new_n992), .B2(G953), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n937), .B1(G898), .B2(new_n224), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT123), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n993), .B(new_n995), .ZN(G69));
  AND2_X1   g810(.A1(new_n857), .A2(new_n719), .ZN(new_n997));
  AND2_X1   g811(.A1(new_n836), .A2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n803), .ZN(new_n999));
  NOR4_X1   g813(.A1(new_n638), .A2(new_n739), .A3(new_n562), .A4(new_n523), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n999), .B1(new_n827), .B2(new_n1000), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n1001), .A2(new_n830), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT126), .ZN(new_n1003));
  NAND4_X1  g817(.A1(new_n998), .A2(new_n1002), .A3(new_n1003), .A4(new_n800), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n836), .A2(new_n1001), .A3(new_n830), .A4(new_n997), .ZN(new_n1005));
  INV_X1    g819(.A(new_n800), .ZN(new_n1006));
  OAI21_X1  g820(.A(KEYINPUT126), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1004), .A2(new_n1007), .A3(new_n224), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n297), .A2(new_n298), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n475), .B1(new_n209), .B2(new_n474), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1008), .B(new_n1011), .C1(new_n688), .C2(new_n224), .ZN(new_n1012));
  INV_X1    g826(.A(new_n374), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n845), .A2(new_n846), .ZN(new_n1014));
  XOR2_X1   g828(.A(new_n1014), .B(KEYINPUT125), .Z(new_n1015));
  NAND4_X1  g829(.A1(new_n1013), .A2(new_n712), .A3(new_n794), .A4(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n836), .A2(new_n830), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n714), .A2(new_n997), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1017), .B1(new_n1018), .B2(KEYINPUT62), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT62), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n714), .A2(KEYINPUT124), .A3(new_n1020), .A4(new_n997), .ZN(new_n1021));
  INV_X1    g835(.A(KEYINPUT124), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1022), .B1(new_n1018), .B2(KEYINPUT62), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1019), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n1024), .A2(new_n224), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1012), .B1(new_n1025), .B2(new_n1011), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n224), .B1(G227), .B2(G900), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1027), .ZN(new_n1029));
  OAI211_X1 g843(.A(new_n1012), .B(new_n1029), .C1(new_n1025), .C2(new_n1011), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1028), .A2(new_n1030), .ZN(G72));
  NAND3_X1  g845(.A1(new_n1004), .A2(new_n1007), .A3(new_n992), .ZN(new_n1032));
  NAND2_X1  g846(.A1(G472), .A2(G902), .ZN(new_n1033));
  XOR2_X1   g847(.A(new_n1033), .B(KEYINPUT63), .Z(new_n1034));
  NAND2_X1  g848(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g849(.A1(new_n1035), .A2(new_n301), .A3(new_n342), .A4(new_n299), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n349), .A2(new_n311), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n873), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1036), .A2(new_n964), .A3(new_n1038), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n1019), .A2(new_n992), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1040));
  INV_X1    g854(.A(KEYINPUT127), .ZN(new_n1041));
  AND3_X1   g855(.A1(new_n1040), .A2(new_n1041), .A3(new_n1034), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1041), .B1(new_n1040), .B2(new_n1034), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n369), .A2(new_n310), .ZN(new_n1044));
  NOR3_X1   g858(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n1039), .A2(new_n1045), .ZN(G57));
endmodule


