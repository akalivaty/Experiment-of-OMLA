

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372,
         n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383,
         n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394,
         n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405,
         n406, n407, n408, n409, n410, n411, n412, n413, n414, n415, n416,
         n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, n427,
         n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438,
         n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
         n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460,
         n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762;

  NOR2_X1 U384 ( .A1(n688), .A2(n687), .ZN(n364) );
  NAND2_X2 U385 ( .A1(n447), .A2(n619), .ZN(n621) );
  XNOR2_X2 U386 ( .A(n428), .B(n427), .ZN(n645) );
  NAND2_X1 U387 ( .A1(n364), .A2(n630), .ZN(n411) );
  XNOR2_X2 U388 ( .A(n508), .B(G469), .ZN(n623) );
  INV_X1 U389 ( .A(KEYINPUT4), .ZN(n461) );
  OR2_X1 U390 ( .A1(n380), .A2(n394), .ZN(n640) );
  NAND2_X1 U391 ( .A1(n453), .A2(n452), .ZN(n654) );
  XNOR2_X1 U392 ( .A(n411), .B(n482), .ZN(n699) );
  XNOR2_X1 U393 ( .A(n588), .B(KEYINPUT38), .ZN(n701) );
  NAND2_X1 U394 ( .A1(n471), .A2(n468), .ZN(n683) );
  XNOR2_X1 U395 ( .A(n738), .B(n465), .ZN(n504) );
  XNOR2_X1 U396 ( .A(n512), .B(n466), .ZN(n465) );
  XNOR2_X1 U397 ( .A(n461), .B(G146), .ZN(n501) );
  XOR2_X1 U398 ( .A(KEYINPUT66), .B(G101), .Z(n512) );
  XNOR2_X1 U399 ( .A(KEYINPUT70), .B(G113), .ZN(n483) );
  INV_X2 U400 ( .A(G953), .ZN(n749) );
  NOR2_X2 U401 ( .A1(n677), .A2(n676), .ZN(n678) );
  NOR2_X1 U402 ( .A1(n668), .A2(n670), .ZN(n704) );
  XNOR2_X1 U403 ( .A(G143), .B(n489), .ZN(n499) );
  XNOR2_X1 U404 ( .A(G128), .B(KEYINPUT80), .ZN(n489) );
  NAND2_X1 U405 ( .A1(n639), .A2(KEYINPUT44), .ZN(n399) );
  AND2_X1 U406 ( .A1(n604), .A2(n442), .ZN(n601) );
  INV_X1 U407 ( .A(KEYINPUT85), .ZN(n442) );
  XNOR2_X1 U408 ( .A(n535), .B(n534), .ZN(n544) );
  XOR2_X1 U409 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n534) );
  XNOR2_X1 U410 ( .A(n533), .B(n532), .ZN(n535) );
  INV_X1 U411 ( .A(KEYINPUT69), .ZN(n532) );
  OR2_X1 U412 ( .A1(G902), .A2(G237), .ZN(n567) );
  XNOR2_X1 U413 ( .A(n431), .B(n494), .ZN(n513) );
  XNOR2_X1 U414 ( .A(n493), .B(n483), .ZN(n431) );
  XNOR2_X1 U415 ( .A(G119), .B(G116), .ZN(n493) );
  XNOR2_X1 U416 ( .A(n443), .B(n540), .ZN(n745) );
  INV_X1 U417 ( .A(G137), .ZN(n502) );
  XNOR2_X1 U418 ( .A(n499), .B(n500), .ZN(n540) );
  INV_X1 U419 ( .A(G134), .ZN(n500) );
  NAND2_X1 U420 ( .A1(n732), .A2(n429), .ZN(n459) );
  NOR2_X1 U421 ( .A1(n646), .A2(n430), .ZN(n429) );
  INV_X1 U422 ( .A(KEYINPUT2), .ZN(n430) );
  XNOR2_X1 U423 ( .A(KEYINPUT84), .B(KEYINPUT2), .ZN(n676) );
  INV_X1 U424 ( .A(KEYINPUT22), .ZN(n620) );
  AND2_X1 U425 ( .A1(n757), .A2(n661), .ZN(n432) );
  XNOR2_X1 U426 ( .A(n381), .B(KEYINPUT67), .ZN(n380) );
  XNOR2_X1 U427 ( .A(n397), .B(n396), .ZN(n395) );
  INV_X1 U428 ( .A(KEYINPUT92), .ZN(n396) );
  AND2_X1 U429 ( .A1(n654), .A2(n365), .ZN(n398) );
  NOR2_X1 U430 ( .A1(n437), .A2(n608), .ZN(n424) );
  XNOR2_X1 U431 ( .A(n385), .B(n583), .ZN(n436) );
  XNOR2_X1 U432 ( .A(KEYINPUT10), .B(n517), .ZN(n747) );
  XOR2_X1 U433 ( .A(KEYINPUT76), .B(G140), .Z(n506) );
  INV_X1 U434 ( .A(KEYINPUT71), .ZN(n466) );
  XNOR2_X1 U435 ( .A(n490), .B(KEYINPUT97), .ZN(n451) );
  XNOR2_X1 U436 ( .A(n480), .B(n479), .ZN(n488) );
  XNOR2_X1 U437 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n479) );
  XNOR2_X1 U438 ( .A(n568), .B(KEYINPUT81), .ZN(n569) );
  XNOR2_X1 U439 ( .A(n592), .B(KEYINPUT19), .ZN(n616) );
  XNOR2_X1 U440 ( .A(n492), .B(G107), .ZN(n738) );
  XNOR2_X1 U441 ( .A(G104), .B(G110), .ZN(n492) );
  XNOR2_X1 U442 ( .A(n513), .B(n495), .ZN(n739) );
  XNOR2_X1 U443 ( .A(KEYINPUT16), .B(G122), .ZN(n495) );
  XNOR2_X1 U444 ( .A(G119), .B(G110), .ZN(n545) );
  XNOR2_X1 U445 ( .A(n417), .B(n373), .ZN(n681) );
  AND2_X1 U446 ( .A1(n387), .A2(n701), .ZN(n417) );
  NOR2_X1 U447 ( .A1(n703), .A2(n388), .ZN(n387) );
  XNOR2_X1 U448 ( .A(n580), .B(KEYINPUT39), .ZN(n610) );
  AND2_X1 U449 ( .A1(n634), .A2(n400), .ZN(n622) );
  NAND2_X1 U450 ( .A1(n470), .A2(n469), .ZN(n468) );
  AND2_X1 U451 ( .A1(n467), .A2(n472), .ZN(n471) );
  NOR2_X1 U452 ( .A1(n362), .A2(G902), .ZN(n469) );
  OR2_X1 U453 ( .A1(n688), .A2(KEYINPUT91), .ZN(n454) );
  XNOR2_X1 U454 ( .A(n444), .B(n745), .ZN(n653) );
  XNOR2_X1 U455 ( .A(n514), .B(n445), .ZN(n444) );
  XNOR2_X1 U456 ( .A(n511), .B(n446), .ZN(n445) );
  XNOR2_X1 U457 ( .A(n539), .B(n425), .ZN(n542) );
  XNOR2_X1 U458 ( .A(n538), .B(n426), .ZN(n425) );
  AND2_X1 U459 ( .A1(n459), .A2(G475), .ZN(n392) );
  AND2_X1 U460 ( .A1(n459), .A2(G469), .ZN(n391) );
  NAND2_X1 U461 ( .A1(n460), .A2(n390), .ZN(n647) );
  AND2_X1 U462 ( .A1(n459), .A2(G210), .ZN(n390) );
  AND2_X1 U463 ( .A1(n384), .A2(n363), .ZN(n383) );
  NAND2_X1 U464 ( .A1(n701), .A2(n700), .ZN(n389) );
  NOR2_X1 U465 ( .A1(n598), .A2(n664), .ZN(n438) );
  XNOR2_X1 U466 ( .A(n481), .B(G125), .ZN(n480) );
  XNOR2_X1 U467 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n481) );
  NAND2_X1 U468 ( .A1(G234), .A2(G237), .ZN(n556) );
  XNOR2_X1 U469 ( .A(KEYINPUT15), .B(G902), .ZN(n565) );
  INV_X1 U470 ( .A(KEYINPUT45), .ZN(n427) );
  NAND2_X1 U471 ( .A1(n640), .A2(n395), .ZN(n428) );
  XOR2_X1 U472 ( .A(G131), .B(G104), .Z(n519) );
  XNOR2_X1 U473 ( .A(n418), .B(G122), .ZN(n518) );
  XNOR2_X1 U474 ( .A(G143), .B(KEYINPUT12), .ZN(n520) );
  XOR2_X1 U475 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n521) );
  NAND2_X1 U476 ( .A1(n412), .A2(n415), .ZN(n646) );
  NOR2_X1 U477 ( .A1(n758), .A2(n416), .ZN(n415) );
  INV_X1 U478 ( .A(n675), .ZN(n416) );
  INV_X1 U479 ( .A(n576), .ZN(n690) );
  INV_X1 U480 ( .A(n700), .ZN(n388) );
  NAND2_X1 U481 ( .A1(n362), .A2(G902), .ZN(n472) );
  XNOR2_X1 U482 ( .A(n512), .B(KEYINPUT75), .ZN(n446) );
  XNOR2_X1 U483 ( .A(G116), .B(G122), .ZN(n536) );
  XOR2_X1 U484 ( .A(KEYINPUT107), .B(G107), .Z(n537) );
  INV_X1 U485 ( .A(KEYINPUT7), .ZN(n426) );
  XNOR2_X1 U486 ( .A(n745), .B(n464), .ZN(n648) );
  XNOR2_X1 U487 ( .A(n504), .B(n507), .ZN(n464) );
  XNOR2_X1 U488 ( .A(n449), .B(n448), .ZN(n566) );
  XNOR2_X1 U489 ( .A(n491), .B(n450), .ZN(n448) );
  XNOR2_X1 U490 ( .A(n739), .B(n496), .ZN(n449) );
  NAND2_X1 U491 ( .A1(n719), .A2(n463), .ZN(n434) );
  AND2_X1 U492 ( .A1(n423), .A2(n624), .ZN(n586) );
  OR2_X1 U493 ( .A1(n575), .A2(n440), .ZN(n604) );
  NAND2_X1 U494 ( .A1(n413), .A2(n441), .ZN(n440) );
  INV_X1 U495 ( .A(n623), .ZN(n441) );
  NOR2_X1 U496 ( .A1(n623), .A2(n687), .ZN(n624) );
  XNOR2_X1 U497 ( .A(n447), .B(KEYINPUT102), .ZN(n379) );
  XNOR2_X1 U498 ( .A(n551), .B(n473), .ZN(n729) );
  XNOR2_X1 U499 ( .A(n548), .B(n547), .ZN(n473) );
  XNOR2_X1 U500 ( .A(n386), .B(KEYINPUT42), .ZN(n760) );
  XNOR2_X1 U501 ( .A(n582), .B(n422), .ZN(n762) );
  INV_X1 U502 ( .A(KEYINPUT40), .ZN(n422) );
  AND2_X1 U503 ( .A1(n610), .A2(n668), .ZN(n582) );
  XNOR2_X1 U504 ( .A(n421), .B(n636), .ZN(n757) );
  NAND2_X1 U505 ( .A1(n634), .A2(n635), .ZN(n421) );
  BUF_X1 U506 ( .A(G113), .Z(n418) );
  NOR2_X1 U507 ( .A1(n600), .A2(n599), .ZN(n670) );
  AND2_X1 U508 ( .A1(n455), .A2(n370), .ZN(n453) );
  NAND2_X1 U509 ( .A1(n410), .A2(n409), .ZN(n407) );
  XNOR2_X1 U510 ( .A(n458), .B(n377), .ZN(n410) );
  XNOR2_X1 U511 ( .A(n724), .B(n414), .ZN(n727) );
  XNOR2_X1 U512 ( .A(n726), .B(n725), .ZN(n414) );
  INV_X1 U513 ( .A(KEYINPUT60), .ZN(n405) );
  NAND2_X1 U514 ( .A1(n408), .A2(n409), .ZN(n406) );
  XNOR2_X1 U515 ( .A(n723), .B(n378), .ZN(n408) );
  INV_X1 U516 ( .A(KEYINPUT122), .ZN(n403) );
  INV_X1 U517 ( .A(KEYINPUT56), .ZN(n401) );
  INV_X1 U518 ( .A(KEYINPUT53), .ZN(n462) );
  XOR2_X1 U519 ( .A(n553), .B(KEYINPUT25), .Z(n362) );
  XNOR2_X1 U520 ( .A(n623), .B(KEYINPUT1), .ZN(n688) );
  AND2_X1 U521 ( .A1(n434), .A2(n749), .ZN(n363) );
  OR2_X1 U522 ( .A1(n628), .A2(n627), .ZN(n365) );
  NOR2_X1 U523 ( .A1(n719), .A2(n463), .ZN(n366) );
  AND2_X1 U524 ( .A1(n459), .A2(G472), .ZN(n367) );
  AND2_X1 U525 ( .A1(n383), .A2(n382), .ZN(n368) );
  NOR2_X1 U526 ( .A1(n576), .A2(n683), .ZN(n369) );
  AND2_X1 U527 ( .A1(n454), .A2(n683), .ZN(n370) );
  XOR2_X1 U528 ( .A(n620), .B(KEYINPUT73), .Z(n371) );
  XOR2_X1 U529 ( .A(KEYINPUT96), .B(n617), .Z(n372) );
  XOR2_X1 U530 ( .A(KEYINPUT41), .B(KEYINPUT110), .Z(n373) );
  XOR2_X1 U531 ( .A(n498), .B(n497), .Z(n374) );
  XOR2_X1 U532 ( .A(n650), .B(n649), .Z(n375) );
  XNOR2_X1 U533 ( .A(KEYINPUT48), .B(KEYINPUT89), .ZN(n376) );
  XOR2_X1 U534 ( .A(n653), .B(n652), .Z(n377) );
  XOR2_X1 U535 ( .A(n722), .B(n721), .Z(n378) );
  INV_X1 U536 ( .A(n731), .ZN(n409) );
  NAND2_X1 U537 ( .A1(n379), .A2(n699), .ZN(n478) );
  NAND2_X1 U538 ( .A1(n379), .A2(n624), .ZN(n625) );
  NOR2_X1 U539 ( .A1(n756), .A2(KEYINPUT44), .ZN(n381) );
  NOR2_X1 U540 ( .A1(n679), .A2(n680), .ZN(n720) );
  NAND2_X1 U541 ( .A1(n679), .A2(n366), .ZN(n382) );
  NAND2_X1 U542 ( .A1(n680), .A2(n366), .ZN(n384) );
  NAND2_X1 U543 ( .A1(n368), .A2(n433), .ZN(n435) );
  NAND2_X1 U544 ( .A1(n760), .A2(n762), .ZN(n385) );
  NAND2_X1 U545 ( .A1(n590), .A2(n681), .ZN(n386) );
  NOR2_X1 U546 ( .A1(n704), .A2(n389), .ZN(n705) );
  AND2_X1 U547 ( .A1(n460), .A2(n459), .ZN(n393) );
  NAND2_X1 U548 ( .A1(n460), .A2(n391), .ZN(n651) );
  NAND2_X1 U549 ( .A1(n460), .A2(n367), .ZN(n458) );
  NAND2_X1 U550 ( .A1(n460), .A2(n392), .ZN(n723) );
  NAND2_X1 U551 ( .A1(n393), .A2(G217), .ZN(n728) );
  NAND2_X1 U552 ( .A1(n393), .A2(G478), .ZN(n724) );
  INV_X1 U553 ( .A(n432), .ZN(n394) );
  NAND2_X1 U554 ( .A1(n399), .A2(n398), .ZN(n397) );
  INV_X1 U555 ( .A(n630), .ZN(n400) );
  AND2_X1 U556 ( .A1(n634), .A2(n369), .ZN(n637) );
  XNOR2_X2 U557 ( .A(n621), .B(n371), .ZN(n634) );
  XNOR2_X1 U558 ( .A(n402), .B(n401), .ZN(G51) );
  NAND2_X1 U559 ( .A1(n419), .A2(n409), .ZN(n402) );
  XNOR2_X1 U560 ( .A(n404), .B(n403), .ZN(G54) );
  NAND2_X1 U561 ( .A1(n420), .A2(n409), .ZN(n404) );
  XNOR2_X1 U562 ( .A(n406), .B(n405), .ZN(G60) );
  XNOR2_X1 U563 ( .A(n407), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X2 U564 ( .A1(n644), .A2(n643), .ZN(n460) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(n443) );
  INV_X1 U566 ( .A(n681), .ZN(n698) );
  XNOR2_X1 U567 ( .A(n609), .B(n376), .ZN(n412) );
  BUF_X1 U568 ( .A(n616), .Z(n413) );
  NOR2_X2 U569 ( .A1(n645), .A2(n748), .ZN(n677) );
  XNOR2_X1 U570 ( .A(n647), .B(n374), .ZN(n419) );
  XNOR2_X1 U571 ( .A(n651), .B(n375), .ZN(n420) );
  NAND2_X1 U572 ( .A1(n729), .A2(n362), .ZN(n467) );
  NOR2_X1 U573 ( .A1(n579), .A2(n578), .ZN(n423) );
  NAND2_X1 U574 ( .A1(n677), .A2(n641), .ZN(n644) );
  NAND2_X1 U575 ( .A1(n424), .A2(n436), .ZN(n609) );
  XNOR2_X1 U576 ( .A(n607), .B(KEYINPUT74), .ZN(n439) );
  NAND2_X1 U577 ( .A1(n638), .A2(n432), .ZN(n639) );
  NAND2_X1 U578 ( .A1(n720), .A2(n463), .ZN(n433) );
  XNOR2_X1 U579 ( .A(n435), .B(n462), .ZN(G75) );
  NAND2_X1 U580 ( .A1(n439), .A2(n438), .ZN(n437) );
  NOR2_X1 U581 ( .A1(n575), .A2(n623), .ZN(n590) );
  INV_X1 U582 ( .A(n604), .ZN(n665) );
  NAND2_X1 U583 ( .A1(n447), .A2(n695), .ZN(n626) );
  XNOR2_X2 U584 ( .A(n474), .B(n372), .ZN(n447) );
  XNOR2_X1 U585 ( .A(n499), .B(n451), .ZN(n450) );
  OR2_X1 U586 ( .A1(n457), .A2(KEYINPUT91), .ZN(n452) );
  NAND2_X1 U587 ( .A1(n457), .A2(n456), .ZN(n455) );
  AND2_X1 U588 ( .A1(n688), .A2(KEYINPUT91), .ZN(n456) );
  XNOR2_X1 U589 ( .A(n622), .B(KEYINPUT90), .ZN(n457) );
  INV_X1 U590 ( .A(n459), .ZN(n680) );
  NOR2_X1 U591 ( .A1(n690), .A2(n573), .ZN(n574) );
  NOR2_X1 U592 ( .A1(n704), .A2(n601), .ZN(n603) );
  INV_X1 U593 ( .A(KEYINPUT119), .ZN(n463) );
  INV_X1 U594 ( .A(n729), .ZN(n470) );
  NAND2_X1 U595 ( .A1(n616), .A2(n615), .ZN(n474) );
  NAND2_X2 U596 ( .A1(n589), .A2(n700), .ZN(n592) );
  XNOR2_X2 U597 ( .A(n475), .B(KEYINPUT35), .ZN(n756) );
  NAND2_X1 U598 ( .A1(n476), .A2(n629), .ZN(n475) );
  XNOR2_X1 U599 ( .A(n478), .B(n477), .ZN(n476) );
  INV_X1 U600 ( .A(KEYINPUT34), .ZN(n477) );
  XNOR2_X1 U601 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n482) );
  INV_X1 U602 ( .A(KEYINPUT59), .ZN(n721) );
  XNOR2_X1 U603 ( .A(n550), .B(n549), .ZN(n551) );
  NOR2_X1 U604 ( .A1(G952), .A2(n749), .ZN(n731) );
  XOR2_X1 U605 ( .A(KEYINPUT95), .B(KEYINPUT94), .Z(n485) );
  XNOR2_X1 U606 ( .A(KEYINPUT55), .B(KEYINPUT83), .ZN(n484) );
  XNOR2_X1 U607 ( .A(n485), .B(n484), .ZN(n486) );
  XOR2_X1 U608 ( .A(n486), .B(KEYINPUT120), .Z(n498) );
  XNOR2_X1 U609 ( .A(n501), .B(KEYINPUT77), .ZN(n487) );
  XNOR2_X1 U610 ( .A(n488), .B(n487), .ZN(n491) );
  NAND2_X1 U611 ( .A1(G224), .A2(n749), .ZN(n490) );
  INV_X1 U612 ( .A(n504), .ZN(n496) );
  XOR2_X1 U613 ( .A(KEYINPUT98), .B(KEYINPUT3), .Z(n494) );
  XNOR2_X1 U614 ( .A(n566), .B(KEYINPUT54), .ZN(n497) );
  INV_X1 U615 ( .A(n565), .ZN(n641) );
  XNOR2_X1 U616 ( .A(n501), .B(G131), .ZN(n503) );
  NAND2_X1 U617 ( .A1(G227), .A2(n749), .ZN(n505) );
  XNOR2_X1 U618 ( .A(n506), .B(n505), .ZN(n507) );
  NOR2_X1 U619 ( .A1(G902), .A2(n648), .ZN(n508) );
  XOR2_X1 U620 ( .A(n623), .B(KEYINPUT1), .Z(n631) );
  NOR2_X1 U621 ( .A1(G953), .A2(G237), .ZN(n524) );
  NAND2_X1 U622 ( .A1(n524), .A2(G210), .ZN(n510) );
  XOR2_X1 U623 ( .A(KEYINPUT103), .B(KEYINPUT5), .Z(n509) );
  XNOR2_X1 U624 ( .A(n510), .B(n509), .ZN(n511) );
  BUF_X1 U625 ( .A(n513), .Z(n514) );
  NOR2_X1 U626 ( .A1(n653), .A2(G902), .ZN(n516) );
  INV_X1 U627 ( .A(G472), .ZN(n515) );
  XNOR2_X2 U628 ( .A(n516), .B(n515), .ZN(n576) );
  XOR2_X1 U629 ( .A(KEYINPUT6), .B(n576), .Z(n630) );
  XOR2_X1 U630 ( .A(G125), .B(G140), .Z(n517) );
  XNOR2_X1 U631 ( .A(G146), .B(n747), .ZN(n550) );
  XNOR2_X1 U632 ( .A(n519), .B(n518), .ZN(n523) );
  XNOR2_X1 U633 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U634 ( .A(n523), .B(n522), .ZN(n528) );
  XOR2_X1 U635 ( .A(KEYINPUT106), .B(KEYINPUT11), .Z(n526) );
  NAND2_X1 U636 ( .A1(n524), .A2(G214), .ZN(n525) );
  XNOR2_X1 U637 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U638 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U639 ( .A(n550), .B(n529), .ZN(n722) );
  NOR2_X1 U640 ( .A1(G902), .A2(n722), .ZN(n531) );
  XNOR2_X1 U641 ( .A(KEYINPUT13), .B(G475), .ZN(n530) );
  XNOR2_X1 U642 ( .A(n531), .B(n530), .ZN(n600) );
  NAND2_X1 U643 ( .A1(G234), .A2(n749), .ZN(n533) );
  NAND2_X1 U644 ( .A1(G217), .A2(n544), .ZN(n539) );
  XNOR2_X1 U645 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U646 ( .A(n540), .B(KEYINPUT9), .ZN(n541) );
  XNOR2_X1 U647 ( .A(n542), .B(n541), .ZN(n726) );
  NOR2_X1 U648 ( .A1(n726), .A2(G902), .ZN(n543) );
  XOR2_X1 U649 ( .A(n543), .B(G478), .Z(n584) );
  INV_X1 U650 ( .A(n584), .ZN(n599) );
  NAND2_X1 U651 ( .A1(n600), .A2(n599), .ZN(n581) );
  NAND2_X1 U652 ( .A1(G221), .A2(n544), .ZN(n548) );
  XOR2_X1 U653 ( .A(G137), .B(G128), .Z(n546) );
  XNOR2_X1 U654 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U655 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n549) );
  NAND2_X1 U656 ( .A1(G234), .A2(n565), .ZN(n552) );
  XNOR2_X1 U657 ( .A(KEYINPUT20), .B(n552), .ZN(n559) );
  NAND2_X1 U658 ( .A1(n559), .A2(G217), .ZN(n553) );
  NOR2_X1 U659 ( .A1(G900), .A2(n749), .ZN(n554) );
  NAND2_X1 U660 ( .A1(n554), .A2(G902), .ZN(n555) );
  NAND2_X1 U661 ( .A1(G952), .A2(n749), .ZN(n612) );
  NAND2_X1 U662 ( .A1(n555), .A2(n612), .ZN(n558) );
  XOR2_X1 U663 ( .A(n556), .B(KEYINPUT14), .Z(n715) );
  INV_X1 U664 ( .A(n715), .ZN(n557) );
  NAND2_X1 U665 ( .A1(n558), .A2(n557), .ZN(n578) );
  NOR2_X1 U666 ( .A1(n683), .A2(n578), .ZN(n561) );
  NAND2_X1 U667 ( .A1(n559), .A2(G221), .ZN(n560) );
  XNOR2_X1 U668 ( .A(KEYINPUT21), .B(n560), .ZN(n618) );
  INV_X1 U669 ( .A(n618), .ZN(n684) );
  NAND2_X1 U670 ( .A1(n561), .A2(n684), .ZN(n573) );
  NOR2_X1 U671 ( .A1(n581), .A2(n573), .ZN(n562) );
  NAND2_X1 U672 ( .A1(n630), .A2(n562), .ZN(n593) );
  NOR2_X1 U673 ( .A1(n631), .A2(n593), .ZN(n563) );
  NAND2_X1 U674 ( .A1(G214), .A2(n567), .ZN(n700) );
  NAND2_X1 U675 ( .A1(n563), .A2(n700), .ZN(n564) );
  XNOR2_X1 U676 ( .A(n564), .B(KEYINPUT43), .ZN(n571) );
  NAND2_X1 U677 ( .A1(n566), .A2(n565), .ZN(n570) );
  NAND2_X1 U678 ( .A1(G210), .A2(n567), .ZN(n568) );
  XNOR2_X2 U679 ( .A(n570), .B(n569), .ZN(n589) );
  INV_X1 U680 ( .A(n589), .ZN(n588) );
  NAND2_X1 U681 ( .A1(n571), .A2(n588), .ZN(n572) );
  XNOR2_X1 U682 ( .A(KEYINPUT109), .B(n572), .ZN(n758) );
  OR2_X1 U683 ( .A1(n584), .A2(n600), .ZN(n703) );
  XOR2_X1 U684 ( .A(KEYINPUT28), .B(n574), .Z(n575) );
  NAND2_X1 U685 ( .A1(n576), .A2(n700), .ZN(n577) );
  XNOR2_X1 U686 ( .A(KEYINPUT30), .B(n577), .ZN(n579) );
  NAND2_X1 U687 ( .A1(n684), .A2(n683), .ZN(n687) );
  NAND2_X1 U688 ( .A1(n586), .A2(n701), .ZN(n580) );
  INV_X1 U689 ( .A(n581), .ZN(n668) );
  XOR2_X1 U690 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n583) );
  NAND2_X1 U691 ( .A1(n584), .A2(n600), .ZN(n585) );
  XOR2_X1 U692 ( .A(KEYINPUT108), .B(n585), .Z(n629) );
  NAND2_X1 U693 ( .A1(n586), .A2(n629), .ZN(n587) );
  NOR2_X1 U694 ( .A1(n588), .A2(n587), .ZN(n664) );
  NAND2_X1 U695 ( .A1(n604), .A2(KEYINPUT47), .ZN(n591) );
  NAND2_X1 U696 ( .A1(n591), .A2(KEYINPUT85), .ZN(n597) );
  NOR2_X1 U697 ( .A1(n593), .A2(n592), .ZN(n595) );
  XOR2_X1 U698 ( .A(KEYINPUT36), .B(KEYINPUT93), .Z(n594) );
  XNOR2_X1 U699 ( .A(n595), .B(n594), .ZN(n596) );
  NAND2_X1 U700 ( .A1(n631), .A2(n596), .ZN(n674) );
  NAND2_X1 U701 ( .A1(n597), .A2(n674), .ZN(n598) );
  INV_X1 U702 ( .A(KEYINPUT47), .ZN(n602) );
  NOR2_X1 U703 ( .A1(n603), .A2(n602), .ZN(n608) );
  XNOR2_X1 U704 ( .A(KEYINPUT86), .B(n704), .ZN(n628) );
  INV_X1 U705 ( .A(n628), .ZN(n606) );
  NOR2_X1 U706 ( .A1(n604), .A2(KEYINPUT47), .ZN(n605) );
  NAND2_X1 U707 ( .A1(n606), .A2(n605), .ZN(n607) );
  NAND2_X1 U708 ( .A1(n610), .A2(n670), .ZN(n675) );
  XNOR2_X1 U709 ( .A(KEYINPUT88), .B(n646), .ZN(n748) );
  NOR2_X1 U710 ( .A1(G898), .A2(n749), .ZN(n611) );
  XOR2_X1 U711 ( .A(KEYINPUT101), .B(n611), .Z(n742) );
  NAND2_X1 U712 ( .A1(n742), .A2(G902), .ZN(n613) );
  AND2_X1 U713 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U714 ( .A1(n614), .A2(n715), .ZN(n615) );
  XOR2_X1 U715 ( .A(KEYINPUT65), .B(KEYINPUT0), .Z(n617) );
  NOR2_X1 U716 ( .A1(n703), .A2(n618), .ZN(n619) );
  NOR2_X1 U717 ( .A1(n576), .A2(n625), .ZN(n657) );
  AND2_X1 U718 ( .A1(n576), .A2(n364), .ZN(n695) );
  XNOR2_X1 U719 ( .A(n626), .B(KEYINPUT31), .ZN(n671) );
  NOR2_X1 U720 ( .A1(n657), .A2(n671), .ZN(n627) );
  INV_X1 U721 ( .A(n756), .ZN(n638) );
  XNOR2_X1 U722 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n636) );
  NOR2_X1 U723 ( .A1(n630), .A2(n683), .ZN(n632) );
  NAND2_X1 U724 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U725 ( .A(n633), .B(KEYINPUT79), .ZN(n635) );
  NAND2_X1 U726 ( .A1(n688), .A2(n637), .ZN(n661) );
  XOR2_X1 U727 ( .A(KEYINPUT87), .B(n641), .Z(n642) );
  NAND2_X1 U728 ( .A1(n642), .A2(KEYINPUT2), .ZN(n643) );
  INV_X1 U729 ( .A(n645), .ZN(n732) );
  XNOR2_X1 U730 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n650) );
  XNOR2_X1 U731 ( .A(n648), .B(KEYINPUT57), .ZN(n649) );
  XOR2_X1 U732 ( .A(KEYINPUT111), .B(KEYINPUT62), .Z(n652) );
  XNOR2_X1 U733 ( .A(G101), .B(n654), .ZN(G3) );
  NAND2_X1 U734 ( .A1(n657), .A2(n668), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n655), .B(KEYINPUT112), .ZN(n656) );
  XNOR2_X1 U736 ( .A(G104), .B(n656), .ZN(G6) );
  XOR2_X1 U737 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n659) );
  NAND2_X1 U738 ( .A1(n657), .A2(n670), .ZN(n658) );
  XNOR2_X1 U739 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U740 ( .A(G107), .B(n660), .ZN(G9) );
  XNOR2_X1 U741 ( .A(G110), .B(n661), .ZN(G12) );
  XOR2_X1 U742 ( .A(G128), .B(KEYINPUT29), .Z(n663) );
  NAND2_X1 U743 ( .A1(n670), .A2(n665), .ZN(n662) );
  XNOR2_X1 U744 ( .A(n663), .B(n662), .ZN(G30) );
  XOR2_X1 U745 ( .A(G143), .B(n664), .Z(G45) );
  XOR2_X1 U746 ( .A(G146), .B(KEYINPUT113), .Z(n667) );
  NAND2_X1 U747 ( .A1(n665), .A2(n668), .ZN(n666) );
  XNOR2_X1 U748 ( .A(n667), .B(n666), .ZN(G48) );
  NAND2_X1 U749 ( .A1(n671), .A2(n668), .ZN(n669) );
  XNOR2_X1 U750 ( .A(n669), .B(n418), .ZN(G15) );
  NAND2_X1 U751 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U752 ( .A(n672), .B(G116), .ZN(G18) );
  XOR2_X1 U753 ( .A(G125), .B(KEYINPUT37), .Z(n673) );
  XNOR2_X1 U754 ( .A(n674), .B(n673), .ZN(G27) );
  XNOR2_X1 U755 ( .A(G134), .B(n675), .ZN(G36) );
  XNOR2_X1 U756 ( .A(n678), .B(KEYINPUT82), .ZN(n679) );
  NAND2_X1 U757 ( .A1(n681), .A2(n699), .ZN(n682) );
  XNOR2_X1 U758 ( .A(n682), .B(KEYINPUT118), .ZN(n718) );
  NOR2_X1 U759 ( .A1(n684), .A2(n683), .ZN(n686) );
  XNOR2_X1 U760 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n685) );
  XNOR2_X1 U761 ( .A(n686), .B(n685), .ZN(n693) );
  NAND2_X1 U762 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U763 ( .A(n689), .B(KEYINPUT50), .ZN(n691) );
  NAND2_X1 U764 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U765 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U766 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U767 ( .A(KEYINPUT51), .B(n696), .Z(n697) );
  NOR2_X1 U768 ( .A1(n698), .A2(n697), .ZN(n711) );
  INV_X1 U769 ( .A(n699), .ZN(n709) );
  NOR2_X1 U770 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U771 ( .A1(n703), .A2(n702), .ZN(n707) );
  XNOR2_X1 U772 ( .A(n705), .B(KEYINPUT116), .ZN(n706) );
  NOR2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n708) );
  NOR2_X1 U774 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U775 ( .A1(n711), .A2(n710), .ZN(n712) );
  XOR2_X1 U776 ( .A(n712), .B(KEYINPUT52), .Z(n713) );
  XNOR2_X1 U777 ( .A(KEYINPUT117), .B(n713), .ZN(n714) );
  NOR2_X1 U778 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U779 ( .A1(n716), .A2(G952), .ZN(n717) );
  NAND2_X1 U780 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U781 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n725) );
  NOR2_X1 U782 ( .A1(n731), .A2(n727), .ZN(G63) );
  XNOR2_X1 U783 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U784 ( .A1(n731), .A2(n730), .ZN(G66) );
  NAND2_X1 U785 ( .A1(n749), .A2(n732), .ZN(n736) );
  NAND2_X1 U786 ( .A1(G953), .A2(G224), .ZN(n733) );
  XNOR2_X1 U787 ( .A(KEYINPUT61), .B(n733), .ZN(n734) );
  NAND2_X1 U788 ( .A1(n734), .A2(G898), .ZN(n735) );
  NAND2_X1 U789 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U790 ( .A(n737), .B(KEYINPUT125), .ZN(n744) );
  XOR2_X1 U791 ( .A(n739), .B(n738), .Z(n740) );
  XNOR2_X1 U792 ( .A(G101), .B(n740), .ZN(n741) );
  NOR2_X1 U793 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U794 ( .A(n744), .B(n743), .Z(G69) );
  XOR2_X1 U795 ( .A(n745), .B(KEYINPUT126), .Z(n746) );
  XNOR2_X1 U796 ( .A(n747), .B(n746), .ZN(n751) );
  XNOR2_X1 U797 ( .A(n751), .B(n748), .ZN(n750) );
  NAND2_X1 U798 ( .A1(n750), .A2(n749), .ZN(n755) );
  XNOR2_X1 U799 ( .A(G227), .B(n751), .ZN(n752) );
  NAND2_X1 U800 ( .A1(n752), .A2(G900), .ZN(n753) );
  NAND2_X1 U801 ( .A1(n753), .A2(G953), .ZN(n754) );
  NAND2_X1 U802 ( .A1(n755), .A2(n754), .ZN(G72) );
  XOR2_X1 U803 ( .A(n756), .B(G122), .Z(G24) );
  XNOR2_X1 U804 ( .A(n757), .B(G119), .ZN(G21) );
  XOR2_X1 U805 ( .A(G140), .B(n758), .Z(n759) );
  XNOR2_X1 U806 ( .A(KEYINPUT114), .B(n759), .ZN(G42) );
  XOR2_X1 U807 ( .A(G137), .B(n760), .Z(n761) );
  XNOR2_X1 U808 ( .A(KEYINPUT127), .B(n761), .ZN(G39) );
  XNOR2_X1 U809 ( .A(G131), .B(n762), .ZN(G33) );
endmodule

