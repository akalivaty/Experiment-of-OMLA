

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778;

  XNOR2_X1 U378 ( .A(n414), .B(n481), .ZN(n413) );
  XNOR2_X1 U379 ( .A(n420), .B(G146), .ZN(n378) );
  BUF_X1 U380 ( .A(n722), .Z(n767) );
  BUF_X1 U381 ( .A(n744), .Z(n750) );
  XOR2_X1 U382 ( .A(n381), .B(n448), .Z(n357) );
  AND2_X1 U383 ( .A1(n472), .A2(n373), .ZN(n358) );
  XNOR2_X2 U384 ( .A(n631), .B(n630), .ZN(n643) );
  INV_X1 U385 ( .A(n572), .ZN(n567) );
  NAND2_X1 U386 ( .A1(n624), .A2(n687), .ZN(n594) );
  INV_X1 U387 ( .A(n624), .ZN(n641) );
  XNOR2_X2 U388 ( .A(n484), .B(n483), .ZN(n485) );
  XOR2_X2 U389 ( .A(G131), .B(G137), .Z(n484) );
  NOR2_X1 U390 ( .A1(n366), .A2(KEYINPUT93), .ZN(n361) );
  NAND2_X1 U391 ( .A1(n422), .A2(n473), .ZN(n366) );
  OR2_X1 U392 ( .A1(n453), .A2(n451), .ZN(n576) );
  NOR2_X1 U393 ( .A1(n452), .A2(n456), .ZN(n451) );
  NOR2_X1 U394 ( .A1(n707), .A2(n357), .ZN(n565) );
  NOR2_X4 U395 ( .A1(n573), .A2(n567), .ZN(n670) );
  AND2_X1 U396 ( .A1(n365), .A2(n364), .ZN(n363) );
  OR2_X1 U397 ( .A1(n453), .A2(n451), .ZN(n380) );
  NOR2_X1 U398 ( .A1(n385), .A2(n432), .ZN(n424) );
  XNOR2_X1 U399 ( .A(n392), .B(KEYINPUT33), .ZN(n717) );
  NOR2_X1 U400 ( .A1(n584), .A2(n396), .ZN(n395) );
  NOR2_X1 U401 ( .A1(n758), .A2(n767), .ZN(n646) );
  NOR2_X1 U402 ( .A1(n722), .A2(n479), .ZN(n478) );
  NAND2_X1 U403 ( .A1(n362), .A2(n361), .ZN(n360) );
  NAND2_X1 U404 ( .A1(n421), .A2(n358), .ZN(n367) );
  NAND2_X1 U405 ( .A1(n460), .A2(n457), .ZN(n456) );
  XNOR2_X1 U406 ( .A(n408), .B(n407), .ZN(n696) );
  XNOR2_X1 U407 ( .A(n600), .B(KEYINPUT6), .ZN(n592) );
  INV_X1 U408 ( .A(n701), .ZN(n589) );
  XNOR2_X1 U409 ( .A(n401), .B(n535), .ZN(n572) );
  XOR2_X1 U410 ( .A(n657), .B(KEYINPUT62), .Z(n659) );
  XNOR2_X1 U411 ( .A(n395), .B(n370), .ZN(n553) );
  XNOR2_X1 U412 ( .A(n480), .B(n486), .ZN(n498) );
  XNOR2_X1 U413 ( .A(n416), .B(G143), .ZN(n499) );
  XNOR2_X1 U414 ( .A(n497), .B(KEYINPUT76), .ZN(n481) );
  XNOR2_X1 U415 ( .A(G128), .B(KEYINPUT4), .ZN(n416) );
  XNOR2_X1 U416 ( .A(G134), .B(KEYINPUT9), .ZN(n528) );
  XOR2_X1 U417 ( .A(G143), .B(G128), .Z(n527) );
  NAND2_X1 U418 ( .A1(n359), .A2(n754), .ZN(n762) );
  XNOR2_X2 U419 ( .A(n504), .B(n359), .ZN(n733) );
  XNOR2_X2 U420 ( .A(n413), .B(n498), .ZN(n359) );
  NAND2_X1 U421 ( .A1(n363), .A2(n360), .ZN(n581) );
  INV_X1 U422 ( .A(n367), .ZN(n362) );
  NAND2_X1 U423 ( .A1(n366), .A2(KEYINPUT93), .ZN(n364) );
  NAND2_X1 U424 ( .A1(n367), .A2(KEYINPUT93), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n527), .B(n526), .ZN(n531) );
  BUF_X1 U426 ( .A(n727), .Z(n368) );
  XNOR2_X2 U427 ( .A(n582), .B(n383), .ZN(n382) );
  XNOR2_X1 U428 ( .A(n548), .B(n442), .ZN(n441) );
  OR2_X2 U429 ( .A1(n741), .A2(G902), .ZN(n443) );
  INV_X1 U430 ( .A(G469), .ZN(n442) );
  OR2_X1 U431 ( .A1(n749), .A2(G902), .ZN(n559) );
  XNOR2_X1 U432 ( .A(G140), .B(KEYINPUT10), .ZN(n410) );
  NAND2_X1 U433 ( .A1(n678), .A2(n400), .ZN(n397) );
  INV_X1 U434 ( .A(KEYINPUT77), .ZN(n400) );
  OR2_X1 U435 ( .A1(n644), .A2(n675), .ZN(n608) );
  INV_X1 U436 ( .A(KEYINPUT111), .ZN(n461) );
  NOR2_X1 U437 ( .A1(G953), .A2(G237), .ZN(n518) );
  XNOR2_X1 U438 ( .A(n405), .B(KEYINPUT89), .ZN(n404) );
  NAND2_X1 U439 ( .A1(n566), .A2(n567), .ZN(n690) );
  XNOR2_X1 U440 ( .A(n440), .B(KEYINPUT34), .ZN(n439) );
  NOR2_X1 U441 ( .A1(n717), .A2(n357), .ZN(n440) );
  INV_X1 U442 ( .A(n615), .ZN(n438) );
  NOR2_X1 U443 ( .A1(n696), .A2(n697), .ZN(n574) );
  OR2_X1 U444 ( .A1(G237), .A2(G902), .ZN(n506) );
  NAND2_X1 U445 ( .A1(n553), .A2(G221), .ZN(n464) );
  XNOR2_X1 U446 ( .A(n429), .B(n763), .ZN(n650) );
  XNOR2_X1 U447 ( .A(n523), .B(n517), .ZN(n429) );
  XNOR2_X1 U448 ( .A(n547), .B(n546), .ZN(n741) );
  XNOR2_X1 U449 ( .A(n417), .B(n499), .ZN(n503) );
  XNOR2_X1 U450 ( .A(n629), .B(KEYINPUT74), .ZN(n630) );
  NAND2_X1 U451 ( .A1(n562), .A2(n433), .ZN(n432) );
  INV_X1 U452 ( .A(n592), .ZN(n433) );
  XNOR2_X1 U453 ( .A(n411), .B(n409), .ZN(n749) );
  XNOR2_X1 U454 ( .A(n464), .B(n412), .ZN(n411) );
  XNOR2_X1 U455 ( .A(n763), .B(n552), .ZN(n409) );
  XNOR2_X1 U456 ( .A(n463), .B(n551), .ZN(n412) );
  XNOR2_X1 U457 ( .A(n533), .B(n402), .ZN(n748) );
  XNOR2_X1 U458 ( .A(n525), .B(KEYINPUT106), .ZN(n533) );
  NAND2_X1 U459 ( .A1(n553), .A2(G217), .ZN(n525) );
  INV_X1 U460 ( .A(G953), .ZN(n507) );
  AND2_X1 U461 ( .A1(n589), .A2(KEYINPUT44), .ZN(n560) );
  AND2_X1 U462 ( .A1(n399), .A2(n398), .ZN(n609) );
  NAND2_X1 U463 ( .A1(n386), .A2(n474), .ZN(n472) );
  NAND2_X1 U464 ( .A1(n668), .A2(n391), .ZN(n577) );
  NOR2_X1 U465 ( .A1(n638), .A2(n461), .ZN(n458) );
  AND2_X1 U466 ( .A1(n459), .A2(n600), .ZN(n457) );
  INV_X1 U467 ( .A(G125), .ZN(n420) );
  XOR2_X1 U468 ( .A(KEYINPUT7), .B(KEYINPUT107), .Z(n529) );
  XOR2_X1 U469 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n520) );
  XOR2_X1 U470 ( .A(KEYINPUT12), .B(G131), .Z(n516) );
  XNOR2_X1 U471 ( .A(G113), .B(G143), .ZN(n515) );
  XNOR2_X1 U472 ( .A(G104), .B(G107), .ZN(n538) );
  XOR2_X1 U473 ( .A(KEYINPUT82), .B(G140), .Z(n539) );
  INV_X1 U474 ( .A(KEYINPUT81), .ZN(n540) );
  XNOR2_X1 U475 ( .A(G101), .B(G110), .ZN(n541) );
  XNOR2_X1 U476 ( .A(n378), .B(n418), .ZN(n417) );
  XNOR2_X1 U477 ( .A(n419), .B(KEYINPUT83), .ZN(n418) );
  INV_X1 U478 ( .A(KEYINPUT95), .ZN(n419) );
  XOR2_X1 U479 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n501) );
  AND2_X1 U480 ( .A1(n574), .A2(n592), .ZN(n392) );
  INV_X1 U481 ( .A(KEYINPUT2), .ZN(n479) );
  INV_X1 U482 ( .A(KEYINPUT0), .ZN(n448) );
  XNOR2_X1 U483 ( .A(n488), .B(G116), .ZN(n447) );
  XNOR2_X1 U484 ( .A(n388), .B(KEYINPUT3), .ZN(n480) );
  XNOR2_X1 U485 ( .A(KEYINPUT73), .B(G119), .ZN(n388) );
  XNOR2_X1 U486 ( .A(G110), .B(KEYINPUT16), .ZN(n497) );
  XNOR2_X1 U487 ( .A(n554), .B(KEYINPUT99), .ZN(n463) );
  XNOR2_X1 U488 ( .A(G119), .B(G137), .ZN(n554) );
  XOR2_X1 U489 ( .A(KEYINPUT24), .B(KEYINPUT100), .Z(n551) );
  INV_X1 U490 ( .A(G234), .ZN(n396) );
  XNOR2_X1 U491 ( .A(n437), .B(n377), .ZN(n578) );
  NAND2_X1 U492 ( .A1(n439), .A2(n438), .ZN(n437) );
  XNOR2_X1 U493 ( .A(KEYINPUT109), .B(G478), .ZN(n535) );
  NOR2_X1 U494 ( .A1(n748), .A2(G902), .ZN(n401) );
  XNOR2_X1 U495 ( .A(n524), .B(n430), .ZN(n566) );
  XNOR2_X1 U496 ( .A(n431), .B(G475), .ZN(n430) );
  INV_X1 U497 ( .A(KEYINPUT13), .ZN(n431) );
  XNOR2_X1 U498 ( .A(n613), .B(n470), .ZN(n469) );
  INV_X1 U499 ( .A(KEYINPUT30), .ZN(n470) );
  INV_X1 U500 ( .A(KEYINPUT67), .ZN(n407) );
  XNOR2_X1 U501 ( .A(n547), .B(n393), .ZN(n657) );
  XNOR2_X1 U502 ( .A(n498), .B(n394), .ZN(n393) );
  XNOR2_X1 U503 ( .A(n447), .B(n487), .ZN(n394) );
  XOR2_X1 U504 ( .A(KEYINPUT103), .B(KEYINPUT5), .Z(n487) );
  XNOR2_X1 U505 ( .A(n650), .B(KEYINPUT59), .ZN(n651) );
  XNOR2_X1 U506 ( .A(n734), .B(KEYINPUT54), .ZN(n735) );
  XOR2_X1 U507 ( .A(KEYINPUT94), .B(n653), .Z(n740) );
  NOR2_X1 U508 ( .A1(n597), .A2(n697), .ZN(n684) );
  NOR2_X1 U509 ( .A1(n572), .A2(n566), .ZN(n675) );
  XNOR2_X1 U510 ( .A(n751), .B(n749), .ZN(n435) );
  XNOR2_X1 U511 ( .A(n747), .B(n748), .ZN(n423) );
  XNOR2_X1 U512 ( .A(n745), .B(n746), .ZN(n434) );
  INV_X1 U513 ( .A(KEYINPUT53), .ZN(n427) );
  INV_X1 U514 ( .A(G119), .ZN(n390) );
  AND2_X1 U515 ( .A1(n536), .A2(n700), .ZN(n369) );
  XNOR2_X1 U516 ( .A(KEYINPUT8), .B(KEYINPUT68), .ZN(n370) );
  OR2_X1 U517 ( .A1(n465), .A2(n696), .ZN(n371) );
  NOR2_X1 U518 ( .A1(n696), .A2(n563), .ZN(n372) );
  NOR2_X1 U519 ( .A1(n563), .A2(n614), .ZN(n468) );
  AND2_X1 U520 ( .A1(n571), .A2(n661), .ZN(n373) );
  AND2_X1 U521 ( .A1(n458), .A2(n462), .ZN(n374) );
  AND2_X1 U522 ( .A1(n560), .A2(n474), .ZN(n375) );
  OR2_X1 U523 ( .A1(KEYINPUT47), .A2(KEYINPUT77), .ZN(n376) );
  INV_X1 U524 ( .A(KEYINPUT66), .ZN(n462) );
  XOR2_X1 U525 ( .A(n575), .B(KEYINPUT88), .Z(n377) );
  XNOR2_X1 U526 ( .A(n378), .B(n410), .ZN(n763) );
  XNOR2_X2 U527 ( .A(n379), .B(n496), .ZN(n414) );
  XNOR2_X2 U528 ( .A(n389), .B(G104), .ZN(n379) );
  XNOR2_X1 U529 ( .A(n379), .B(KEYINPUT11), .ZN(n522) );
  XNOR2_X1 U530 ( .A(G122), .B(KEYINPUT108), .ZN(n526) );
  NAND2_X1 U531 ( .A1(n604), .A2(n514), .ZN(n381) );
  NAND2_X1 U532 ( .A1(n604), .A2(n514), .ZN(n449) );
  XNOR2_X1 U533 ( .A(n532), .B(n534), .ZN(n402) );
  XNOR2_X1 U534 ( .A(n449), .B(n448), .ZN(n471) );
  AND2_X1 U535 ( .A1(n469), .A2(n688), .ZN(n444) );
  INV_X1 U536 ( .A(n382), .ZN(n758) );
  XOR2_X1 U537 ( .A(KEYINPUT87), .B(KEYINPUT45), .Z(n383) );
  NAND2_X1 U538 ( .A1(n380), .A2(n375), .ZN(n473) );
  NOR2_X1 U539 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X2 U540 ( .A(n628), .B(KEYINPUT42), .ZN(n778) );
  NOR2_X2 U541 ( .A1(n691), .A2(n690), .ZN(n626) );
  BUF_X1 U542 ( .A(n476), .Z(n384) );
  XNOR2_X1 U543 ( .A(n537), .B(KEYINPUT22), .ZN(n385) );
  XNOR2_X1 U544 ( .A(n424), .B(KEYINPUT32), .ZN(n476) );
  XNOR2_X1 U545 ( .A(n537), .B(KEYINPUT22), .ZN(n561) );
  AND2_X1 U546 ( .A1(n387), .A2(KEYINPUT65), .ZN(n475) );
  NAND2_X1 U547 ( .A1(n454), .A2(n455), .ZN(n453) );
  NAND2_X1 U548 ( .A1(n476), .A2(KEYINPUT44), .ZN(n387) );
  INV_X1 U549 ( .A(n387), .ZN(n386) );
  INV_X2 U550 ( .A(G122), .ZN(n389) );
  XNOR2_X1 U551 ( .A(n384), .B(n390), .ZN(n775) );
  INV_X1 U552 ( .A(n384), .ZN(n391) );
  INV_X1 U553 ( .A(n584), .ZN(n768) );
  OR2_X1 U554 ( .A1(n644), .A2(n397), .ZN(n399) );
  INV_X1 U555 ( .A(n608), .ZN(n692) );
  NAND2_X1 U556 ( .A1(n608), .A2(n376), .ZN(n398) );
  NAND2_X1 U557 ( .A1(n778), .A2(n403), .ZN(n445) );
  XNOR2_X1 U558 ( .A(n403), .B(G131), .ZN(G33) );
  XNOR2_X2 U559 ( .A(n446), .B(KEYINPUT40), .ZN(n403) );
  NAND2_X1 U560 ( .A1(n404), .A2(n777), .ZN(n722) );
  NAND2_X1 U561 ( .A1(n406), .A2(n686), .ZN(n405) );
  XNOR2_X1 U562 ( .A(n426), .B(n636), .ZN(n406) );
  NOR2_X1 U563 ( .A1(n696), .A2(n467), .ZN(n466) );
  NAND2_X1 U564 ( .A1(n701), .A2(n700), .ZN(n408) );
  XNOR2_X2 U565 ( .A(n559), .B(n558), .ZN(n701) );
  NAND2_X1 U566 ( .A1(n450), .A2(n458), .ZN(n415) );
  NAND2_X1 U567 ( .A1(n450), .A2(n374), .ZN(n455) );
  NAND2_X1 U568 ( .A1(n415), .A2(KEYINPUT66), .ZN(n452) );
  NAND2_X1 U569 ( .A1(n578), .A2(KEYINPUT44), .ZN(n421) );
  XNOR2_X1 U570 ( .A(n425), .B(KEYINPUT79), .ZN(n727) );
  NAND2_X1 U571 ( .A1(n477), .A2(n475), .ZN(n422) );
  NOR2_X2 U572 ( .A1(n635), .A2(n684), .ZN(n426) );
  NOR2_X1 U573 ( .A1(n423), .A2(n752), .ZN(G63) );
  NAND2_X1 U574 ( .A1(n382), .A2(n478), .ZN(n425) );
  NAND2_X1 U575 ( .A1(n561), .A2(n461), .ZN(n460) );
  NAND2_X1 U576 ( .A1(n744), .A2(G210), .ZN(n736) );
  AND2_X2 U577 ( .A1(n649), .A2(n648), .ZN(n744) );
  NAND2_X1 U578 ( .A1(n456), .A2(n462), .ZN(n454) );
  OR2_X2 U579 ( .A1(n627), .A2(n718), .ZN(n628) );
  XNOR2_X1 U580 ( .A(n445), .B(n632), .ZN(n633) );
  XNOR2_X2 U581 ( .A(n625), .B(n641), .ZN(n688) );
  XNOR2_X1 U582 ( .A(n428), .B(n427), .ZN(G75) );
  NAND2_X1 U583 ( .A1(n732), .A2(n507), .ZN(n428) );
  NOR2_X1 U584 ( .A1(n434), .A2(n752), .ZN(G54) );
  NOR2_X1 U585 ( .A1(n435), .A2(n752), .ZN(G66) );
  NAND2_X1 U586 ( .A1(n471), .A2(n369), .ZN(n537) );
  XNOR2_X2 U587 ( .A(n505), .B(n482), .ZN(n624) );
  NAND2_X1 U588 ( .A1(n436), .A2(n740), .ZN(n660) );
  XNOR2_X1 U589 ( .A(n658), .B(n659), .ZN(n436) );
  XNOR2_X2 U590 ( .A(n443), .B(n441), .ZN(n602) );
  NAND2_X1 U591 ( .A1(n466), .A2(n444), .ZN(n631) );
  NAND2_X1 U592 ( .A1(n643), .A2(n675), .ZN(n446) );
  XNOR2_X2 U593 ( .A(n764), .B(G146), .ZN(n547) );
  XNOR2_X2 U594 ( .A(n594), .B(KEYINPUT19), .ZN(n604) );
  INV_X1 U595 ( .A(n561), .ZN(n450) );
  NOR2_X1 U596 ( .A1(n385), .A2(n638), .ZN(n570) );
  NAND2_X1 U597 ( .A1(n638), .A2(n461), .ZN(n459) );
  NOR2_X2 U598 ( .A1(n733), .A2(n648), .ZN(n505) );
  XNOR2_X2 U599 ( .A(n499), .B(n485), .ZN(n764) );
  NAND2_X1 U600 ( .A1(n468), .A2(n469), .ZN(n465) );
  INV_X1 U601 ( .A(n468), .ZN(n467) );
  XNOR2_X2 U602 ( .A(G953), .B(KEYINPUT64), .ZN(n584) );
  NAND2_X1 U603 ( .A1(n576), .A2(n560), .ZN(n477) );
  INV_X1 U604 ( .A(KEYINPUT65), .ZN(n474) );
  XNOR2_X1 U605 ( .A(n736), .B(n735), .ZN(n737) );
  NAND2_X1 U606 ( .A1(G210), .A2(n506), .ZN(n482) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(n542) );
  INV_X1 U608 ( .A(KEYINPUT35), .ZN(n575) );
  INV_X1 U609 ( .A(n604), .ZN(n605) );
  XNOR2_X1 U610 ( .A(n652), .B(n651), .ZN(n654) );
  XNOR2_X1 U611 ( .A(G134), .B(KEYINPUT69), .ZN(n483) );
  XNOR2_X1 U612 ( .A(G113), .B(G101), .ZN(n486) );
  AND2_X1 U613 ( .A1(n518), .A2(G210), .ZN(n488) );
  NOR2_X1 U614 ( .A1(G902), .A2(n657), .ZN(n490) );
  XNOR2_X1 U615 ( .A(KEYINPUT75), .B(G472), .ZN(n489) );
  XNOR2_X1 U616 ( .A(n490), .B(n489), .ZN(n612) );
  INV_X1 U617 ( .A(n612), .ZN(n600) );
  INV_X1 U618 ( .A(n600), .ZN(n704) );
  XOR2_X1 U619 ( .A(KEYINPUT102), .B(KEYINPUT21), .Z(n494) );
  XOR2_X2 U620 ( .A(G902), .B(KEYINPUT15), .Z(n648) );
  INV_X1 U621 ( .A(n648), .ZN(n491) );
  NAND2_X1 U622 ( .A1(G234), .A2(n491), .ZN(n492) );
  XNOR2_X1 U623 ( .A(KEYINPUT20), .B(n492), .ZN(n555) );
  NAND2_X1 U624 ( .A1(n555), .A2(G221), .ZN(n493) );
  XNOR2_X1 U625 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U626 ( .A(KEYINPUT101), .B(n495), .Z(n700) );
  INV_X1 U627 ( .A(n700), .ZN(n588) );
  XNOR2_X2 U628 ( .A(G116), .B(G107), .ZN(n534) );
  INV_X1 U629 ( .A(n534), .ZN(n496) );
  NAND2_X1 U630 ( .A1(G224), .A2(n768), .ZN(n500) );
  XNOR2_X1 U631 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U632 ( .A(n503), .B(n502), .ZN(n504) );
  NAND2_X1 U633 ( .A1(G214), .A2(n506), .ZN(n687) );
  NOR2_X1 U634 ( .A1(G898), .A2(n507), .ZN(n753) );
  NAND2_X1 U635 ( .A1(G234), .A2(G237), .ZN(n508) );
  XNOR2_X1 U636 ( .A(n508), .B(KEYINPUT14), .ZN(n510) );
  NAND2_X1 U637 ( .A1(n510), .A2(G902), .ZN(n509) );
  XNOR2_X1 U638 ( .A(n509), .B(KEYINPUT97), .ZN(n583) );
  NAND2_X1 U639 ( .A1(n753), .A2(n583), .ZN(n513) );
  NAND2_X1 U640 ( .A1(G952), .A2(n510), .ZN(n511) );
  XNOR2_X1 U641 ( .A(n511), .B(KEYINPUT96), .ZN(n715) );
  NOR2_X1 U642 ( .A1(G953), .A2(n715), .ZN(n587) );
  INV_X1 U643 ( .A(n587), .ZN(n512) );
  NAND2_X1 U644 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U645 ( .A(n516), .B(n515), .ZN(n517) );
  NAND2_X1 U646 ( .A1(n518), .A2(G214), .ZN(n519) );
  XNOR2_X1 U647 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U648 ( .A(n522), .B(n521), .ZN(n523) );
  NOR2_X1 U649 ( .A1(G902), .A2(n650), .ZN(n524) );
  XNOR2_X1 U650 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U651 ( .A(n531), .B(n530), .Z(n532) );
  INV_X1 U652 ( .A(n690), .ZN(n536) );
  NAND2_X1 U653 ( .A1(G227), .A2(n768), .ZN(n545) );
  XNOR2_X1 U654 ( .A(n539), .B(n538), .ZN(n543) );
  XNOR2_X1 U655 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U656 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U657 ( .A(KEYINPUT71), .B(KEYINPUT72), .ZN(n548) );
  XOR2_X2 U658 ( .A(KEYINPUT1), .B(n602), .Z(n697) );
  INV_X1 U659 ( .A(n697), .ZN(n638) );
  XOR2_X1 U660 ( .A(KEYINPUT23), .B(KEYINPUT98), .Z(n550) );
  XNOR2_X1 U661 ( .A(G110), .B(G128), .ZN(n549) );
  XNOR2_X1 U662 ( .A(n550), .B(n549), .ZN(n552) );
  XOR2_X1 U663 ( .A(KEYINPUT25), .B(KEYINPUT80), .Z(n557) );
  NAND2_X1 U664 ( .A1(n555), .A2(G217), .ZN(n556) );
  XNOR2_X1 U665 ( .A(n557), .B(n556), .ZN(n558) );
  NOR2_X1 U666 ( .A1(n697), .A2(n701), .ZN(n562) );
  INV_X1 U667 ( .A(n602), .ZN(n563) );
  NOR2_X1 U668 ( .A1(n704), .A2(n357), .ZN(n564) );
  NAND2_X1 U669 ( .A1(n372), .A2(n564), .ZN(n664) );
  NAND2_X1 U670 ( .A1(n704), .A2(n574), .ZN(n707) );
  XNOR2_X1 U671 ( .A(n565), .B(KEYINPUT31), .ZN(n680) );
  NAND2_X1 U672 ( .A1(n664), .A2(n680), .ZN(n568) );
  INV_X1 U673 ( .A(n566), .ZN(n573) );
  XNOR2_X1 U674 ( .A(KEYINPUT110), .B(n670), .ZN(n644) );
  NAND2_X1 U675 ( .A1(n568), .A2(n608), .ZN(n571) );
  NOR2_X1 U676 ( .A1(n592), .A2(n589), .ZN(n569) );
  NAND2_X1 U677 ( .A1(n570), .A2(n569), .ZN(n661) );
  NAND2_X1 U678 ( .A1(n573), .A2(n572), .ZN(n615) );
  NAND2_X1 U679 ( .A1(n380), .A2(n589), .ZN(n668) );
  NOR2_X1 U680 ( .A1(KEYINPUT44), .A2(n577), .ZN(n579) );
  INV_X1 U681 ( .A(n578), .ZN(n776) );
  NAND2_X1 U682 ( .A1(n579), .A2(n776), .ZN(n580) );
  NAND2_X1 U683 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U684 ( .A(KEYINPUT70), .B(KEYINPUT48), .ZN(n636) );
  INV_X1 U685 ( .A(n675), .ZN(n678) );
  NAND2_X1 U686 ( .A1(n584), .A2(n583), .ZN(n585) );
  NOR2_X1 U687 ( .A1(G900), .A2(n585), .ZN(n586) );
  NOR2_X1 U688 ( .A1(n587), .A2(n586), .ZN(n614) );
  NOR2_X1 U689 ( .A1(n614), .A2(n588), .ZN(n590) );
  NAND2_X1 U690 ( .A1(n590), .A2(n589), .ZN(n599) );
  NOR2_X1 U691 ( .A1(n678), .A2(n599), .ZN(n591) );
  NAND2_X1 U692 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U693 ( .A(KEYINPUT112), .B(n593), .ZN(n637) );
  NOR2_X1 U694 ( .A1(n637), .A2(n594), .ZN(n596) );
  XNOR2_X1 U695 ( .A(KEYINPUT113), .B(KEYINPUT36), .ZN(n595) );
  XNOR2_X1 U696 ( .A(n596), .B(n595), .ZN(n597) );
  INV_X1 U697 ( .A(KEYINPUT84), .ZN(n619) );
  NOR2_X1 U698 ( .A1(n608), .A2(n619), .ZN(n598) );
  NOR2_X1 U699 ( .A1(KEYINPUT77), .A2(n598), .ZN(n606) );
  NOR2_X1 U700 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U701 ( .A(n601), .B(KEYINPUT28), .ZN(n603) );
  NAND2_X1 U702 ( .A1(n603), .A2(n602), .ZN(n627) );
  NOR2_X1 U703 ( .A1(n627), .A2(n605), .ZN(n676) );
  NAND2_X1 U704 ( .A1(n606), .A2(n676), .ZN(n607) );
  NAND2_X1 U705 ( .A1(n607), .A2(KEYINPUT47), .ZN(n611) );
  NAND2_X1 U706 ( .A1(n609), .A2(n676), .ZN(n610) );
  AND2_X1 U707 ( .A1(n611), .A2(n610), .ZN(n623) );
  NAND2_X1 U708 ( .A1(n612), .A2(n687), .ZN(n613) );
  NOR2_X1 U709 ( .A1(n371), .A2(n615), .ZN(n616) );
  NAND2_X1 U710 ( .A1(n624), .A2(n616), .ZN(n674) );
  NAND2_X1 U711 ( .A1(n692), .A2(KEYINPUT47), .ZN(n617) );
  NAND2_X1 U712 ( .A1(n674), .A2(n617), .ZN(n618) );
  NAND2_X1 U713 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U714 ( .A1(n674), .A2(KEYINPUT84), .ZN(n620) );
  NAND2_X1 U715 ( .A1(n621), .A2(n620), .ZN(n622) );
  AND2_X1 U716 ( .A1(n623), .A2(n622), .ZN(n634) );
  XNOR2_X1 U717 ( .A(KEYINPUT38), .B(KEYINPUT78), .ZN(n625) );
  NAND2_X1 U718 ( .A1(n688), .A2(n687), .ZN(n691) );
  XNOR2_X1 U719 ( .A(KEYINPUT41), .B(n626), .ZN(n718) );
  XNOR2_X1 U720 ( .A(KEYINPUT92), .B(KEYINPUT39), .ZN(n629) );
  XNOR2_X1 U721 ( .A(KEYINPUT46), .B(KEYINPUT91), .ZN(n632) );
  NAND2_X1 U722 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U723 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U724 ( .A1(n639), .A2(n687), .ZN(n640) );
  XNOR2_X1 U725 ( .A(n640), .B(KEYINPUT43), .ZN(n642) );
  NAND2_X1 U726 ( .A1(n642), .A2(n641), .ZN(n686) );
  NAND2_X1 U727 ( .A1(n643), .A2(n644), .ZN(n645) );
  XNOR2_X1 U728 ( .A(KEYINPUT114), .B(n645), .ZN(n777) );
  NOR2_X1 U729 ( .A1(n646), .A2(KEYINPUT2), .ZN(n647) );
  NOR2_X1 U730 ( .A1(n727), .A2(n647), .ZN(n649) );
  NAND2_X1 U731 ( .A1(n744), .A2(G475), .ZN(n652) );
  NOR2_X1 U732 ( .A1(n768), .A2(G952), .ZN(n653) );
  NAND2_X1 U733 ( .A1(n654), .A2(n740), .ZN(n656) );
  INV_X1 U734 ( .A(KEYINPUT60), .ZN(n655) );
  XNOR2_X1 U735 ( .A(n656), .B(n655), .ZN(G60) );
  NAND2_X1 U736 ( .A1(n744), .A2(G472), .ZN(n658) );
  XNOR2_X1 U737 ( .A(n660), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U738 ( .A(G101), .B(n661), .ZN(G3) );
  NOR2_X1 U739 ( .A1(n678), .A2(n664), .ZN(n663) );
  XNOR2_X1 U740 ( .A(G104), .B(KEYINPUT115), .ZN(n662) );
  XNOR2_X1 U741 ( .A(n663), .B(n662), .ZN(G6) );
  INV_X1 U742 ( .A(n670), .ZN(n681) );
  NOR2_X1 U743 ( .A1(n681), .A2(n664), .ZN(n666) );
  XNOR2_X1 U744 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n665) );
  XNOR2_X1 U745 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U746 ( .A(G107), .B(n667), .ZN(G9) );
  XNOR2_X1 U747 ( .A(G110), .B(KEYINPUT116), .ZN(n669) );
  XNOR2_X1 U748 ( .A(n669), .B(n668), .ZN(G12) );
  XOR2_X1 U749 ( .A(G128), .B(KEYINPUT29), .Z(n672) );
  NAND2_X1 U750 ( .A1(n676), .A2(n670), .ZN(n671) );
  XNOR2_X1 U751 ( .A(n672), .B(n671), .ZN(G30) );
  XOR2_X1 U752 ( .A(G143), .B(KEYINPUT117), .Z(n673) );
  XNOR2_X1 U753 ( .A(n674), .B(n673), .ZN(G45) );
  NAND2_X1 U754 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U755 ( .A(n677), .B(G146), .ZN(G48) );
  NOR2_X1 U756 ( .A1(n678), .A2(n680), .ZN(n679) );
  XOR2_X1 U757 ( .A(G113), .B(n679), .Z(G15) );
  NOR2_X1 U758 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U759 ( .A(KEYINPUT118), .B(n682), .Z(n683) );
  XNOR2_X1 U760 ( .A(G116), .B(n683), .ZN(G18) );
  XNOR2_X1 U761 ( .A(n684), .B(G125), .ZN(n685) );
  XNOR2_X1 U762 ( .A(n685), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U763 ( .A(G140), .B(n686), .ZN(G42) );
  NOR2_X1 U764 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U765 ( .A1(n690), .A2(n689), .ZN(n694) );
  NOR2_X1 U766 ( .A1(n692), .A2(n691), .ZN(n693) );
  NOR2_X1 U767 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U768 ( .A1(n717), .A2(n695), .ZN(n712) );
  AND2_X1 U769 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U770 ( .A(n698), .B(KEYINPUT50), .ZN(n699) );
  XNOR2_X1 U771 ( .A(n699), .B(KEYINPUT119), .ZN(n706) );
  NOR2_X1 U772 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U773 ( .A(KEYINPUT49), .B(n702), .Z(n703) );
  NOR2_X1 U774 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U775 ( .A1(n706), .A2(n705), .ZN(n708) );
  NAND2_X1 U776 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U777 ( .A(KEYINPUT51), .B(n709), .ZN(n710) );
  NOR2_X1 U778 ( .A1(n710), .A2(n718), .ZN(n711) );
  NOR2_X1 U779 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U780 ( .A(n713), .B(KEYINPUT52), .ZN(n714) );
  NOR2_X1 U781 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U782 ( .A(n716), .B(KEYINPUT120), .ZN(n720) );
  NOR2_X1 U783 ( .A1(n718), .A2(n717), .ZN(n719) );
  NOR2_X1 U784 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U785 ( .A(n721), .B(KEYINPUT121), .ZN(n730) );
  XNOR2_X1 U786 ( .A(KEYINPUT2), .B(KEYINPUT85), .ZN(n724) );
  NAND2_X1 U787 ( .A1(n767), .A2(n724), .ZN(n723) );
  XNOR2_X1 U788 ( .A(n723), .B(KEYINPUT86), .ZN(n726) );
  NAND2_X1 U789 ( .A1(n724), .A2(n758), .ZN(n725) );
  NAND2_X1 U790 ( .A1(n726), .A2(n725), .ZN(n728) );
  NOR2_X1 U791 ( .A1(n728), .A2(n368), .ZN(n729) );
  XNOR2_X1 U792 ( .A(n731), .B(KEYINPUT122), .ZN(n732) );
  XNOR2_X1 U793 ( .A(n733), .B(KEYINPUT55), .ZN(n734) );
  NAND2_X1 U794 ( .A1(n737), .A2(n740), .ZN(n739) );
  XOR2_X1 U795 ( .A(KEYINPUT90), .B(KEYINPUT56), .Z(n738) );
  XNOR2_X1 U796 ( .A(n739), .B(n738), .ZN(G51) );
  INV_X1 U797 ( .A(n740), .ZN(n752) );
  XNOR2_X1 U798 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n743) );
  XNOR2_X1 U799 ( .A(n741), .B(KEYINPUT57), .ZN(n742) );
  XNOR2_X1 U800 ( .A(n743), .B(n742), .ZN(n746) );
  NAND2_X1 U801 ( .A1(n750), .A2(G469), .ZN(n745) );
  NAND2_X1 U802 ( .A1(G478), .A2(n750), .ZN(n747) );
  NAND2_X1 U803 ( .A1(G217), .A2(n750), .ZN(n751) );
  INV_X1 U804 ( .A(n753), .ZN(n754) );
  NAND2_X1 U805 ( .A1(G953), .A2(G224), .ZN(n755) );
  XNOR2_X1 U806 ( .A(KEYINPUT61), .B(n755), .ZN(n756) );
  NAND2_X1 U807 ( .A1(n756), .A2(G898), .ZN(n757) );
  XOR2_X1 U808 ( .A(KEYINPUT124), .B(n757), .Z(n760) );
  NOR2_X1 U809 ( .A1(G953), .A2(n758), .ZN(n759) );
  NOR2_X1 U810 ( .A1(n760), .A2(n759), .ZN(n761) );
  XNOR2_X1 U811 ( .A(n762), .B(n761), .ZN(G69) );
  XNOR2_X1 U812 ( .A(n764), .B(n763), .ZN(n770) );
  INV_X1 U813 ( .A(n770), .ZN(n765) );
  XNOR2_X1 U814 ( .A(KEYINPUT125), .B(n765), .ZN(n766) );
  XNOR2_X1 U815 ( .A(n767), .B(n766), .ZN(n769) );
  NAND2_X1 U816 ( .A1(n769), .A2(n768), .ZN(n774) );
  XNOR2_X1 U817 ( .A(G227), .B(n770), .ZN(n771) );
  NAND2_X1 U818 ( .A1(n771), .A2(G900), .ZN(n772) );
  NAND2_X1 U819 ( .A1(n772), .A2(G953), .ZN(n773) );
  NAND2_X1 U820 ( .A1(n774), .A2(n773), .ZN(G72) );
  XNOR2_X1 U821 ( .A(n775), .B(KEYINPUT126), .ZN(G21) );
  XNOR2_X1 U822 ( .A(G122), .B(n776), .ZN(G24) );
  XNOR2_X1 U823 ( .A(G134), .B(n777), .ZN(G36) );
  XNOR2_X1 U824 ( .A(G137), .B(n778), .ZN(G39) );
endmodule

