

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786;

  INV_X1 U377 ( .A(n680), .ZN(n355) );
  OR2_X1 U378 ( .A1(n662), .A2(n663), .ZN(n435) );
  NAND2_X1 U379 ( .A1(n586), .A2(n563), .ZN(n694) );
  OR2_X1 U380 ( .A1(n742), .A2(G902), .ZN(n512) );
  XNOR2_X1 U381 ( .A(n356), .B(n355), .ZN(G51) );
  NAND2_X1 U382 ( .A1(n381), .A2(n378), .ZN(n356) );
  AND2_X1 U383 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U384 ( .A1(n580), .A2(n368), .ZN(n590) );
  BUF_X1 U385 ( .A(n741), .Z(n752) );
  NAND2_X1 U386 ( .A1(n448), .A2(n447), .ZN(n589) );
  AND2_X2 U387 ( .A1(n386), .A2(KEYINPUT64), .ZN(n385) );
  AND2_X2 U388 ( .A1(n638), .A2(n637), .ZN(n383) );
  NAND2_X2 U389 ( .A1(n436), .A2(n459), .ZN(n421) );
  XNOR2_X2 U390 ( .A(n512), .B(n511), .ZN(n655) );
  NOR2_X1 U391 ( .A1(n724), .A2(n723), .ZN(n382) );
  AND2_X1 U392 ( .A1(n390), .A2(n389), .ZN(n388) );
  AND2_X1 U393 ( .A1(n647), .A2(n781), .ZN(n665) );
  XNOR2_X1 U394 ( .A(n633), .B(KEYINPUT42), .ZN(n786) );
  AND2_X1 U395 ( .A1(n439), .A2(n440), .ZN(n418) );
  NAND2_X1 U396 ( .A1(n450), .A2(n449), .ZN(n447) );
  XNOR2_X1 U397 ( .A(n382), .B(n631), .ZN(n734) );
  NOR2_X1 U398 ( .A1(n628), .A2(n627), .ZN(n629) );
  XNOR2_X1 U399 ( .A(n651), .B(n443), .ZN(n460) );
  XNOR2_X1 U400 ( .A(n627), .B(n531), .ZN(n570) );
  NAND2_X1 U401 ( .A1(n428), .A2(n398), .ZN(n627) );
  XNOR2_X1 U402 ( .A(n364), .B(n476), .ZN(n580) );
  AND2_X1 U403 ( .A1(n425), .A2(n399), .ZN(n398) );
  XNOR2_X1 U404 ( .A(n528), .B(n763), .ZN(n677) );
  INV_X1 U405 ( .A(n668), .ZN(n357) );
  XNOR2_X1 U406 ( .A(G128), .B(KEYINPUT97), .ZN(n463) );
  XNOR2_X1 U407 ( .A(n359), .B(n360), .ZN(G60) );
  NAND2_X1 U408 ( .A1(n379), .A2(n378), .ZN(n359) );
  XNOR2_X1 U409 ( .A(KEYINPUT123), .B(KEYINPUT60), .ZN(n360) );
  XNOR2_X1 U410 ( .A(n361), .B(n362), .ZN(G57) );
  NAND2_X1 U411 ( .A1(n380), .A2(n378), .ZN(n361) );
  XNOR2_X1 U412 ( .A(KEYINPUT92), .B(KEYINPUT63), .ZN(n362) );
  XNOR2_X2 U413 ( .A(KEYINPUT69), .B(G131), .ZN(n542) );
  XNOR2_X1 U414 ( .A(n515), .B(KEYINPUT10), .ZN(n769) );
  XNOR2_X2 U415 ( .A(n583), .B(n582), .ZN(n733) );
  NOR2_X1 U416 ( .A1(n599), .A2(n598), .ZN(n602) );
  NOR2_X1 U417 ( .A1(n725), .A2(KEYINPUT47), .ZN(n619) );
  INV_X1 U418 ( .A(G237), .ZN(n492) );
  XNOR2_X1 U419 ( .A(n411), .B(n410), .ZN(n409) );
  INV_X1 U420 ( .A(KEYINPUT48), .ZN(n410) );
  INV_X1 U421 ( .A(KEYINPUT38), .ZN(n397) );
  NOR2_X1 U422 ( .A1(n428), .A2(n397), .ZN(n396) );
  XNOR2_X1 U423 ( .A(n498), .B(G472), .ZN(n499) );
  XNOR2_X1 U424 ( .A(G146), .B(G125), .ZN(n515) );
  XNOR2_X1 U425 ( .A(KEYINPUT18), .B(KEYINPUT94), .ZN(n517) );
  XNOR2_X1 U426 ( .A(KEYINPUT83), .B(KEYINPUT17), .ZN(n518) );
  XNOR2_X1 U427 ( .A(n516), .B(n515), .ZN(n415) );
  XNOR2_X1 U428 ( .A(n419), .B(KEYINPUT73), .ZN(n516) );
  NAND2_X1 U429 ( .A1(n514), .A2(G224), .ZN(n419) );
  INV_X1 U430 ( .A(G953), .ZN(n514) );
  OR2_X2 U431 ( .A1(n677), .A2(n426), .ZN(n425) );
  NAND2_X1 U432 ( .A1(n427), .A2(n357), .ZN(n426) );
  INV_X1 U433 ( .A(n529), .ZN(n427) );
  XNOR2_X1 U434 ( .A(G116), .B(G107), .ZN(n556) );
  AND2_X1 U435 ( .A1(n445), .A2(n610), .ZN(n444) );
  XNOR2_X1 U436 ( .A(KEYINPUT67), .B(KEYINPUT19), .ZN(n531) );
  INV_X1 U437 ( .A(KEYINPUT22), .ZN(n454) );
  NAND2_X1 U438 ( .A1(n725), .A2(KEYINPUT47), .ZN(n611) );
  AND2_X1 U439 ( .A1(n611), .A2(n438), .ZN(n437) );
  INV_X1 U440 ( .A(KEYINPUT85), .ZN(n438) );
  XNOR2_X1 U441 ( .A(n636), .B(n371), .ZN(n637) );
  INV_X1 U442 ( .A(KEYINPUT76), .ZN(n412) );
  XNOR2_X1 U443 ( .A(n493), .B(KEYINPUT81), .ZN(n537) );
  NAND2_X1 U444 ( .A1(n668), .A2(KEYINPUT2), .ZN(n406) );
  XNOR2_X1 U445 ( .A(G143), .B(G140), .ZN(n533) );
  XNOR2_X1 U446 ( .A(n542), .B(G134), .ZN(n502) );
  XNOR2_X1 U447 ( .A(G137), .B(G140), .ZN(n501) );
  INV_X1 U448 ( .A(n701), .ZN(n387) );
  NAND2_X1 U449 ( .A1(G234), .A2(G237), .ZN(n480) );
  XOR2_X1 U450 ( .A(KEYINPUT79), .B(KEYINPUT14), .Z(n481) );
  INV_X1 U451 ( .A(KEYINPUT108), .ZN(n443) );
  AND2_X1 U452 ( .A1(n694), .A2(n697), .ZN(n725) );
  AND2_X1 U453 ( .A1(n409), .A2(n363), .ZN(n402) );
  AND2_X1 U454 ( .A1(n434), .A2(n435), .ZN(n420) );
  AND2_X1 U455 ( .A1(n662), .A2(n663), .ZN(n433) );
  NAND2_X1 U456 ( .A1(n394), .A2(n392), .ZN(n721) );
  NOR2_X1 U457 ( .A1(n396), .A2(n395), .ZN(n394) );
  XNOR2_X1 U458 ( .A(n655), .B(KEYINPUT1), .ZN(n581) );
  OR2_X2 U459 ( .A1(n581), .A2(n706), .ZN(n651) );
  XOR2_X1 U460 ( .A(n600), .B(KEYINPUT30), .Z(n601) );
  INV_X1 U461 ( .A(G902), .ZN(n559) );
  XNOR2_X1 U462 ( .A(KEYINPUT72), .B(KEYINPUT3), .ZN(n525) );
  XNOR2_X1 U463 ( .A(n453), .B(n452), .ZN(n524) );
  INV_X1 U464 ( .A(G104), .ZN(n452) );
  XNOR2_X1 U465 ( .A(G122), .B(G113), .ZN(n453) );
  XNOR2_X1 U466 ( .A(KEYINPUT23), .B(KEYINPUT96), .ZN(n467) );
  XNOR2_X1 U467 ( .A(n502), .B(n501), .ZN(n772) );
  XNOR2_X1 U468 ( .A(n520), .B(n404), .ZN(n528) );
  XNOR2_X1 U469 ( .A(n415), .B(n519), .ZN(n520) );
  XNOR2_X1 U470 ( .A(n594), .B(n593), .ZN(n628) );
  NOR2_X1 U471 ( .A1(n654), .A2(n370), .ZN(n449) );
  NOR2_X2 U472 ( .A1(n570), .A2(n569), .ZN(n571) );
  INV_X2 U473 ( .A(G953), .ZN(n774) );
  XNOR2_X1 U474 ( .A(n555), .B(n422), .ZN(n748) );
  XNOR2_X1 U475 ( .A(n554), .B(n558), .ZN(n422) );
  NOR2_X1 U476 ( .A1(n773), .A2(n405), .ZN(n704) );
  NAND2_X1 U477 ( .A1(n579), .A2(n580), .ZN(n647) );
  AND2_X1 U478 ( .A1(n640), .A2(KEYINPUT2), .ZN(n363) );
  AND2_X1 U479 ( .A1(n753), .A2(n559), .ZN(n364) );
  NOR2_X1 U480 ( .A1(n575), .A2(n712), .ZN(n365) );
  NOR2_X1 U481 ( .A1(n728), .A2(n733), .ZN(n366) );
  AND2_X1 U482 ( .A1(n610), .A2(KEYINPUT85), .ZN(n367) );
  AND2_X1 U483 ( .A1(n486), .A2(n603), .ZN(n368) );
  INV_X1 U484 ( .A(n598), .ZN(n399) );
  NOR2_X1 U485 ( .A1(n574), .A2(n592), .ZN(n369) );
  XOR2_X1 U486 ( .A(n585), .B(KEYINPUT34), .Z(n370) );
  XOR2_X1 U487 ( .A(KEYINPUT90), .B(KEYINPUT46), .Z(n371) );
  XOR2_X1 U488 ( .A(n682), .B(KEYINPUT59), .Z(n372) );
  XOR2_X1 U489 ( .A(n677), .B(n676), .Z(n373) );
  XOR2_X1 U490 ( .A(n684), .B(n685), .Z(n374) );
  AND2_X1 U491 ( .A1(n406), .A2(n673), .ZN(n375) );
  AND2_X1 U492 ( .A1(KEYINPUT91), .A2(KEYINPUT44), .ZN(n376) );
  AND2_X1 U493 ( .A1(n679), .A2(G953), .ZN(n757) );
  INV_X1 U494 ( .A(n757), .ZN(n378) );
  NAND2_X1 U495 ( .A1(n377), .A2(n383), .ZN(n411) );
  XNOR2_X1 U496 ( .A(n626), .B(n412), .ZN(n377) );
  XNOR2_X1 U497 ( .A(n683), .B(n372), .ZN(n379) );
  XNOR2_X1 U498 ( .A(n686), .B(n374), .ZN(n380) );
  XNOR2_X1 U499 ( .A(n678), .B(n373), .ZN(n381) );
  NAND2_X1 U500 ( .A1(n385), .A2(n387), .ZN(n384) );
  BUF_X4 U501 ( .A(n599), .Z(n650) );
  AND2_X1 U502 ( .A1(n446), .A2(n444), .ZN(n448) );
  NAND2_X2 U503 ( .A1(n388), .A2(n384), .ZN(n741) );
  NAND2_X1 U504 ( .A1(n687), .A2(n437), .ZN(n417) );
  NAND2_X1 U505 ( .A1(n408), .A2(n407), .ZN(n391) );
  NAND2_X1 U506 ( .A1(n391), .A2(n406), .ZN(n386) );
  NAND2_X1 U507 ( .A1(n391), .A2(n375), .ZN(n389) );
  NAND2_X1 U508 ( .A1(n701), .A2(n673), .ZN(n390) );
  XNOR2_X2 U509 ( .A(n672), .B(n671), .ZN(n701) );
  NAND2_X1 U510 ( .A1(n428), .A2(n425), .ZN(n607) );
  NAND2_X1 U511 ( .A1(n428), .A2(n393), .ZN(n392) );
  AND2_X1 U512 ( .A1(n425), .A2(n397), .ZN(n393) );
  NOR2_X1 U513 ( .A1(n425), .A2(n397), .ZN(n395) );
  INV_X1 U514 ( .A(n400), .ZN(n405) );
  AND2_X1 U515 ( .A1(n400), .A2(n668), .ZN(n407) );
  XNOR2_X2 U516 ( .A(n421), .B(KEYINPUT45), .ZN(n400) );
  NAND2_X1 U517 ( .A1(n400), .A2(n670), .ZN(n672) );
  NAND2_X1 U518 ( .A1(n400), .A2(n774), .ZN(n761) );
  NAND2_X1 U519 ( .A1(n409), .A2(n640), .ZN(n669) );
  XNOR2_X1 U520 ( .A(n402), .B(n401), .ZN(n670) );
  INV_X1 U521 ( .A(KEYINPUT89), .ZN(n401) );
  NAND2_X1 U522 ( .A1(n403), .A2(n423), .ZN(n635) );
  NAND2_X1 U523 ( .A1(n403), .A2(n424), .ZN(n699) );
  XNOR2_X2 U524 ( .A(n634), .B(KEYINPUT39), .ZN(n403) );
  XNOR2_X1 U525 ( .A(n404), .B(G146), .ZN(n508) );
  XNOR2_X2 U526 ( .A(n768), .B(G101), .ZN(n404) );
  XNOR2_X1 U527 ( .A(n702), .B(n442), .ZN(n408) );
  NAND2_X1 U528 ( .A1(n413), .A2(n367), .ZN(n439) );
  NAND2_X1 U529 ( .A1(n413), .A2(n610), .ZN(n687) );
  XNOR2_X2 U530 ( .A(n609), .B(KEYINPUT113), .ZN(n413) );
  XNOR2_X2 U531 ( .A(n414), .B(KEYINPUT115), .ZN(n782) );
  NAND2_X1 U532 ( .A1(n630), .A2(n575), .ZN(n414) );
  OR2_X2 U533 ( .A1(n651), .A2(n650), .ZN(n653) );
  XNOR2_X1 U534 ( .A(n416), .B(KEYINPUT31), .ZN(n696) );
  NOR2_X1 U535 ( .A1(n716), .A2(n654), .ZN(n416) );
  NAND2_X1 U536 ( .A1(n620), .A2(KEYINPUT47), .ZN(n613) );
  AND2_X1 U537 ( .A1(n430), .A2(n429), .ZN(n428) );
  NAND2_X1 U538 ( .A1(n433), .A2(n432), .ZN(n431) );
  NAND2_X1 U539 ( .A1(n418), .A2(n417), .ZN(n615) );
  NAND2_X1 U540 ( .A1(n451), .A2(n608), .ZN(n609) );
  AND2_X2 U541 ( .A1(n606), .A2(n605), .ZN(n451) );
  XNOR2_X1 U542 ( .A(n457), .B(KEYINPUT28), .ZN(n456) );
  NAND2_X1 U543 ( .A1(n420), .A2(n431), .ZN(n436) );
  AND2_X2 U544 ( .A1(n456), .A2(n513), .ZN(n632) );
  INV_X1 U545 ( .A(n694), .ZN(n423) );
  INV_X1 U546 ( .A(n697), .ZN(n424) );
  NAND2_X1 U547 ( .A1(n529), .A2(n668), .ZN(n429) );
  NAND2_X1 U548 ( .A1(n677), .A2(n529), .ZN(n430) );
  NAND2_X1 U549 ( .A1(n649), .A2(KEYINPUT44), .ZN(n432) );
  NAND2_X1 U550 ( .A1(n649), .A2(n376), .ZN(n434) );
  NAND2_X1 U551 ( .A1(n441), .A2(KEYINPUT85), .ZN(n440) );
  INV_X1 U552 ( .A(n611), .ZN(n441) );
  INV_X1 U553 ( .A(KEYINPUT80), .ZN(n442) );
  XNOR2_X2 U554 ( .A(n669), .B(KEYINPUT88), .ZN(n702) );
  NAND2_X1 U555 ( .A1(n654), .A2(n370), .ZN(n445) );
  NAND2_X1 U556 ( .A1(n733), .A2(n370), .ZN(n446) );
  INV_X1 U557 ( .A(n733), .ZN(n450) );
  NAND2_X1 U558 ( .A1(n451), .A2(n721), .ZN(n634) );
  INV_X1 U559 ( .A(n580), .ZN(n641) );
  INV_X1 U560 ( .A(n524), .ZN(n535) );
  NAND2_X1 U561 ( .A1(n576), .A2(n369), .ZN(n660) );
  XNOR2_X2 U562 ( .A(n573), .B(n454), .ZN(n576) );
  XNOR2_X1 U563 ( .A(n455), .B(G119), .ZN(n489) );
  XNOR2_X2 U564 ( .A(G116), .B(KEYINPUT99), .ZN(n455) );
  NAND2_X2 U565 ( .A1(n632), .A2(n532), .ZN(n620) );
  NOR2_X2 U566 ( .A1(n650), .A2(n590), .ZN(n457) );
  NOR2_X1 U567 ( .A1(n642), .A2(n592), .ZN(n458) );
  OR2_X1 U568 ( .A1(n667), .A2(n666), .ZN(n459) );
  INV_X1 U569 ( .A(KEYINPUT78), .ZN(n618) );
  NAND2_X1 U570 ( .A1(n774), .A2(n492), .ZN(n493) );
  OR2_X2 U571 ( .A1(n684), .A2(G902), .ZN(n500) );
  XOR2_X1 U572 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n462) );
  NAND2_X1 U573 ( .A1(G234), .A2(n774), .ZN(n461) );
  XNOR2_X1 U574 ( .A(n462), .B(n461), .ZN(n550) );
  NAND2_X1 U575 ( .A1(n550), .A2(G221), .ZN(n466) );
  XNOR2_X1 U576 ( .A(n463), .B(KEYINPUT24), .ZN(n464) );
  XNOR2_X1 U577 ( .A(n464), .B(n501), .ZN(n465) );
  XNOR2_X1 U578 ( .A(n466), .B(n465), .ZN(n470) );
  XNOR2_X2 U579 ( .A(G119), .B(G110), .ZN(n522) );
  XNOR2_X1 U580 ( .A(n522), .B(n467), .ZN(n468) );
  XNOR2_X1 U581 ( .A(n769), .B(n468), .ZN(n469) );
  XNOR2_X1 U582 ( .A(n470), .B(n469), .ZN(n753) );
  INV_X1 U583 ( .A(KEYINPUT15), .ZN(n471) );
  XNOR2_X1 U584 ( .A(n471), .B(G902), .ZN(n668) );
  NAND2_X1 U585 ( .A1(n357), .A2(G234), .ZN(n473) );
  INV_X1 U586 ( .A(KEYINPUT20), .ZN(n472) );
  XNOR2_X1 U587 ( .A(n473), .B(n472), .ZN(n478) );
  INV_X1 U588 ( .A(n478), .ZN(n474) );
  AND2_X1 U589 ( .A1(n474), .A2(G217), .ZN(n475) );
  XNOR2_X1 U590 ( .A(n475), .B(KEYINPUT25), .ZN(n476) );
  INV_X1 U591 ( .A(G221), .ZN(n477) );
  OR2_X1 U592 ( .A1(n478), .A2(n477), .ZN(n479) );
  XNOR2_X1 U593 ( .A(n479), .B(KEYINPUT21), .ZN(n710) );
  INV_X1 U594 ( .A(n710), .ZN(n486) );
  XNOR2_X1 U595 ( .A(n481), .B(n480), .ZN(n484) );
  NAND2_X1 U596 ( .A1(G902), .A2(n484), .ZN(n565) );
  NOR2_X1 U597 ( .A1(G900), .A2(n565), .ZN(n482) );
  NAND2_X1 U598 ( .A1(G953), .A2(n482), .ZN(n483) );
  XNOR2_X1 U599 ( .A(n483), .B(KEYINPUT110), .ZN(n485) );
  NAND2_X1 U600 ( .A1(G952), .A2(n484), .ZN(n732) );
  OR2_X1 U601 ( .A1(n732), .A2(G953), .ZN(n566) );
  NAND2_X1 U602 ( .A1(n485), .A2(n566), .ZN(n603) );
  XNOR2_X2 U603 ( .A(G113), .B(G137), .ZN(n488) );
  XNOR2_X2 U604 ( .A(KEYINPUT5), .B(KEYINPUT98), .ZN(n487) );
  XNOR2_X1 U605 ( .A(n488), .B(n487), .ZN(n490) );
  XNOR2_X1 U606 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U607 ( .A(n491), .B(n502), .ZN(n496) );
  NAND2_X1 U608 ( .A1(n537), .A2(G210), .ZN(n494) );
  XNOR2_X1 U609 ( .A(n494), .B(n525), .ZN(n495) );
  XNOR2_X1 U610 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X2 U611 ( .A(G143), .B(G128), .ZN(n552) );
  XNOR2_X2 U612 ( .A(n552), .B(KEYINPUT4), .ZN(n768) );
  XNOR2_X1 U613 ( .A(n497), .B(n508), .ZN(n684) );
  INV_X1 U614 ( .A(KEYINPUT100), .ZN(n498) );
  XNOR2_X2 U615 ( .A(n500), .B(n499), .ZN(n599) );
  NAND2_X1 U616 ( .A1(G227), .A2(n774), .ZN(n503) );
  XNOR2_X1 U617 ( .A(n503), .B(G104), .ZN(n506) );
  XOR2_X1 U618 ( .A(KEYINPUT73), .B(G107), .Z(n504) );
  XNOR2_X1 U619 ( .A(G110), .B(n504), .ZN(n505) );
  XNOR2_X1 U620 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U621 ( .A(n772), .B(n507), .ZN(n509) );
  XNOR2_X1 U622 ( .A(n508), .B(n509), .ZN(n742) );
  XNOR2_X1 U623 ( .A(KEYINPUT71), .B(G469), .ZN(n510) );
  XNOR2_X1 U624 ( .A(n510), .B(KEYINPUT70), .ZN(n511) );
  INV_X1 U625 ( .A(n655), .ZN(n513) );
  XNOR2_X1 U626 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U627 ( .A(KEYINPUT75), .B(KEYINPUT16), .ZN(n521) );
  XNOR2_X1 U628 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U629 ( .A(n523), .B(n524), .ZN(n527) );
  XNOR2_X1 U630 ( .A(n556), .B(n525), .ZN(n526) );
  XNOR2_X1 U631 ( .A(n527), .B(n526), .ZN(n763) );
  NAND2_X1 U632 ( .A1(n559), .A2(n492), .ZN(n530) );
  NAND2_X1 U633 ( .A1(n530), .A2(G210), .ZN(n529) );
  AND2_X1 U634 ( .A1(n530), .A2(G214), .ZN(n598) );
  INV_X1 U635 ( .A(n570), .ZN(n532) );
  XOR2_X1 U636 ( .A(KEYINPUT102), .B(KEYINPUT11), .Z(n534) );
  XNOR2_X1 U637 ( .A(n534), .B(n533), .ZN(n536) );
  XNOR2_X1 U638 ( .A(n536), .B(n535), .ZN(n541) );
  XOR2_X1 U639 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n539) );
  NAND2_X1 U640 ( .A1(n537), .A2(G214), .ZN(n538) );
  XNOR2_X1 U641 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U642 ( .A(n541), .B(n540), .ZN(n545) );
  XNOR2_X1 U643 ( .A(n542), .B(KEYINPUT104), .ZN(n543) );
  XNOR2_X1 U644 ( .A(n769), .B(n543), .ZN(n544) );
  XNOR2_X1 U645 ( .A(n545), .B(n544), .ZN(n682) );
  NAND2_X1 U646 ( .A1(n682), .A2(n559), .ZN(n549) );
  XOR2_X1 U647 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n547) );
  XNOR2_X1 U648 ( .A(KEYINPUT13), .B(G475), .ZN(n546) );
  XOR2_X1 U649 ( .A(n547), .B(n546), .Z(n548) );
  XNOR2_X1 U650 ( .A(n549), .B(n548), .ZN(n586) );
  NAND2_X1 U651 ( .A1(G217), .A2(n550), .ZN(n551) );
  XNOR2_X1 U652 ( .A(G134), .B(n551), .ZN(n555) );
  XNOR2_X1 U653 ( .A(G122), .B(KEYINPUT107), .ZN(n553) );
  XNOR2_X1 U654 ( .A(n552), .B(n553), .ZN(n554) );
  XNOR2_X1 U655 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n557) );
  XNOR2_X1 U656 ( .A(n557), .B(n556), .ZN(n558) );
  NAND2_X1 U657 ( .A1(n748), .A2(n559), .ZN(n560) );
  XNOR2_X1 U658 ( .A(n560), .B(G478), .ZN(n587) );
  INV_X1 U659 ( .A(n587), .ZN(n563) );
  OR2_X1 U660 ( .A1(n586), .A2(n563), .ZN(n697) );
  NOR2_X1 U661 ( .A1(n620), .A2(n697), .ZN(n562) );
  XNOR2_X1 U662 ( .A(G128), .B(KEYINPUT29), .ZN(n561) );
  XNOR2_X1 U663 ( .A(n562), .B(n561), .ZN(G30) );
  NOR2_X1 U664 ( .A1(n620), .A2(n694), .ZN(n564) );
  XOR2_X1 U665 ( .A(G146), .B(n564), .Z(G48) );
  OR2_X1 U666 ( .A1(n774), .A2(G898), .ZN(n764) );
  OR2_X1 U667 ( .A1(n764), .A2(n565), .ZN(n567) );
  NAND2_X1 U668 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U669 ( .A(n568), .B(KEYINPUT95), .ZN(n569) );
  XNOR2_X2 U670 ( .A(n571), .B(KEYINPUT0), .ZN(n584) );
  OR2_X1 U671 ( .A1(n586), .A2(n587), .ZN(n723) );
  NOR2_X1 U672 ( .A1(n723), .A2(n710), .ZN(n572) );
  NAND2_X1 U673 ( .A1(n584), .A2(n572), .ZN(n573) );
  INV_X1 U674 ( .A(n581), .ZN(n575) );
  INV_X1 U675 ( .A(n575), .ZN(n707) );
  NAND2_X1 U676 ( .A1(n707), .A2(n641), .ZN(n574) );
  XNOR2_X2 U677 ( .A(n650), .B(KEYINPUT6), .ZN(n592) );
  XNOR2_X1 U678 ( .A(n660), .B(G101), .ZN(G3) );
  INV_X1 U679 ( .A(n650), .ZN(n712) );
  NAND2_X1 U680 ( .A1(n576), .A2(n365), .ZN(n578) );
  INV_X1 U681 ( .A(KEYINPUT66), .ZN(n577) );
  XNOR2_X1 U682 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U683 ( .A(n647), .B(G110), .ZN(G12) );
  OR2_X1 U684 ( .A1(n580), .A2(n710), .ZN(n706) );
  NAND2_X1 U685 ( .A1(n460), .A2(n592), .ZN(n583) );
  XNOR2_X1 U686 ( .A(KEYINPUT109), .B(KEYINPUT33), .ZN(n582) );
  INV_X1 U687 ( .A(n584), .ZN(n654) );
  INV_X1 U688 ( .A(KEYINPUT74), .ZN(n585) );
  AND2_X1 U689 ( .A1(n587), .A2(n586), .ZN(n610) );
  INV_X1 U690 ( .A(KEYINPUT35), .ZN(n588) );
  XNOR2_X2 U691 ( .A(n589), .B(n588), .ZN(n648) );
  XNOR2_X1 U692 ( .A(n648), .B(G122), .ZN(G24) );
  NOR2_X1 U693 ( .A1(n694), .A2(n590), .ZN(n591) );
  NAND2_X1 U694 ( .A1(n592), .A2(n591), .ZN(n594) );
  INV_X1 U695 ( .A(KEYINPUT111), .ZN(n593) );
  NAND2_X1 U696 ( .A1(n707), .A2(n399), .ZN(n595) );
  OR2_X1 U697 ( .A1(n628), .A2(n595), .ZN(n596) );
  XNOR2_X1 U698 ( .A(n596), .B(KEYINPUT43), .ZN(n597) );
  NAND2_X1 U699 ( .A1(n597), .A2(n607), .ZN(n639) );
  XNOR2_X1 U700 ( .A(n639), .B(G140), .ZN(G42) );
  INV_X1 U701 ( .A(KEYINPUT112), .ZN(n600) );
  XNOR2_X1 U702 ( .A(n602), .B(n601), .ZN(n606) );
  NAND2_X1 U703 ( .A1(n513), .A2(n603), .ZN(n604) );
  NOR2_X1 U704 ( .A1(n604), .A2(n706), .ZN(n605) );
  INV_X1 U705 ( .A(n607), .ZN(n608) );
  INV_X1 U706 ( .A(KEYINPUT87), .ZN(n612) );
  XNOR2_X1 U707 ( .A(n613), .B(n612), .ZN(n614) );
  NAND2_X1 U708 ( .A1(n615), .A2(n614), .ZN(n617) );
  INV_X1 U709 ( .A(KEYINPUT86), .ZN(n616) );
  XNOR2_X1 U710 ( .A(n617), .B(n616), .ZN(n625) );
  XNOR2_X1 U711 ( .A(n619), .B(n618), .ZN(n621) );
  NOR2_X1 U712 ( .A1(n621), .A2(n620), .ZN(n623) );
  INV_X1 U713 ( .A(KEYINPUT77), .ZN(n622) );
  XOR2_X1 U714 ( .A(n623), .B(n622), .Z(n624) );
  NAND2_X1 U715 ( .A1(n625), .A2(n624), .ZN(n626) );
  XNOR2_X1 U716 ( .A(n629), .B(KEYINPUT36), .ZN(n630) );
  INV_X1 U717 ( .A(n782), .ZN(n638) );
  NAND2_X1 U718 ( .A1(n721), .A2(n399), .ZN(n724) );
  XOR2_X1 U719 ( .A(KEYINPUT41), .B(KEYINPUT114), .Z(n631) );
  NAND2_X1 U720 ( .A1(n734), .A2(n632), .ZN(n633) );
  XNOR2_X1 U721 ( .A(n635), .B(KEYINPUT40), .ZN(n785) );
  NAND2_X1 U722 ( .A1(n786), .A2(n785), .ZN(n636) );
  AND2_X1 U723 ( .A1(n639), .A2(n699), .ZN(n640) );
  OR2_X1 U724 ( .A1(n707), .A2(n641), .ZN(n642) );
  NAND2_X1 U725 ( .A1(n576), .A2(n458), .ZN(n646) );
  XNOR2_X1 U726 ( .A(KEYINPUT84), .B(KEYINPUT32), .ZN(n644) );
  INV_X1 U727 ( .A(KEYINPUT65), .ZN(n643) );
  XNOR2_X1 U728 ( .A(n644), .B(n643), .ZN(n645) );
  XNOR2_X1 U729 ( .A(n646), .B(n645), .ZN(n781) );
  NAND2_X1 U730 ( .A1(n665), .A2(n648), .ZN(n649) );
  INV_X1 U731 ( .A(KEYINPUT101), .ZN(n652) );
  XNOR2_X1 U732 ( .A(n653), .B(n652), .ZN(n716) );
  OR2_X1 U733 ( .A1(n706), .A2(n655), .ZN(n656) );
  NOR2_X1 U734 ( .A1(n712), .A2(n656), .ZN(n657) );
  NAND2_X1 U735 ( .A1(n584), .A2(n657), .ZN(n689) );
  NAND2_X1 U736 ( .A1(n696), .A2(n689), .ZN(n659) );
  INV_X1 U737 ( .A(n725), .ZN(n658) );
  NAND2_X1 U738 ( .A1(n659), .A2(n658), .ZN(n661) );
  INV_X1 U739 ( .A(KEYINPUT91), .ZN(n663) );
  INV_X1 U740 ( .A(n648), .ZN(n667) );
  INV_X1 U741 ( .A(KEYINPUT44), .ZN(n664) );
  NAND2_X1 U742 ( .A1(n665), .A2(n664), .ZN(n666) );
  INV_X1 U743 ( .A(KEYINPUT82), .ZN(n671) );
  INV_X1 U744 ( .A(KEYINPUT64), .ZN(n673) );
  NAND2_X1 U745 ( .A1(n741), .A2(G210), .ZN(n678) );
  XOR2_X1 U746 ( .A(KEYINPUT93), .B(KEYINPUT55), .Z(n675) );
  XNOR2_X1 U747 ( .A(KEYINPUT54), .B(KEYINPUT120), .ZN(n674) );
  XOR2_X1 U748 ( .A(n675), .B(n674), .Z(n676) );
  INV_X1 U749 ( .A(G952), .ZN(n679) );
  XOR2_X1 U750 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n680) );
  NAND2_X1 U751 ( .A1(n741), .A2(G475), .ZN(n683) );
  NAND2_X1 U752 ( .A1(n741), .A2(G472), .ZN(n686) );
  XNOR2_X1 U753 ( .A(KEYINPUT116), .B(KEYINPUT62), .ZN(n685) );
  XNOR2_X1 U754 ( .A(n687), .B(G143), .ZN(G45) );
  NOR2_X1 U755 ( .A1(n689), .A2(n694), .ZN(n688) );
  XOR2_X1 U756 ( .A(G104), .B(n688), .Z(G6) );
  NOR2_X1 U757 ( .A1(n689), .A2(n697), .ZN(n693) );
  XOR2_X1 U758 ( .A(KEYINPUT117), .B(KEYINPUT27), .Z(n691) );
  XNOR2_X1 U759 ( .A(G107), .B(KEYINPUT26), .ZN(n690) );
  XNOR2_X1 U760 ( .A(n691), .B(n690), .ZN(n692) );
  XNOR2_X1 U761 ( .A(n693), .B(n692), .ZN(G9) );
  NOR2_X1 U762 ( .A1(n694), .A2(n696), .ZN(n695) );
  XOR2_X1 U763 ( .A(G113), .B(n695), .Z(G15) );
  NOR2_X1 U764 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U765 ( .A(G116), .B(n698), .Z(G18) );
  INV_X1 U766 ( .A(n699), .ZN(n700) );
  XOR2_X1 U767 ( .A(G134), .B(n700), .Z(G36) );
  INV_X1 U768 ( .A(n702), .ZN(n703) );
  INV_X1 U769 ( .A(n703), .ZN(n773) );
  NOR2_X1 U770 ( .A1(n704), .A2(KEYINPUT2), .ZN(n705) );
  NOR2_X1 U771 ( .A1(n701), .A2(n705), .ZN(n738) );
  INV_X1 U772 ( .A(n734), .ZN(n720) );
  NAND2_X1 U773 ( .A1(n707), .A2(n706), .ZN(n709) );
  XOR2_X1 U774 ( .A(KEYINPUT119), .B(KEYINPUT50), .Z(n708) );
  XNOR2_X1 U775 ( .A(n709), .B(n708), .ZN(n715) );
  NAND2_X1 U776 ( .A1(n580), .A2(n710), .ZN(n711) );
  XNOR2_X1 U777 ( .A(n711), .B(KEYINPUT49), .ZN(n713) );
  NOR2_X1 U778 ( .A1(n713), .A2(n712), .ZN(n714) );
  NAND2_X1 U779 ( .A1(n715), .A2(n714), .ZN(n717) );
  NAND2_X1 U780 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U781 ( .A(KEYINPUT51), .B(n718), .ZN(n719) );
  NOR2_X1 U782 ( .A1(n720), .A2(n719), .ZN(n729) );
  NOR2_X1 U783 ( .A1(n721), .A2(n399), .ZN(n722) );
  NOR2_X1 U784 ( .A1(n723), .A2(n722), .ZN(n727) );
  NOR2_X1 U785 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U786 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U787 ( .A1(n729), .A2(n366), .ZN(n730) );
  XNOR2_X1 U788 ( .A(n730), .B(KEYINPUT52), .ZN(n731) );
  NOR2_X1 U789 ( .A1(n732), .A2(n731), .ZN(n736) );
  AND2_X1 U790 ( .A1(n734), .A2(n450), .ZN(n735) );
  OR2_X1 U791 ( .A1(n736), .A2(n735), .ZN(n737) );
  OR2_X1 U792 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U793 ( .A1(n739), .A2(G953), .ZN(n740) );
  XNOR2_X1 U794 ( .A(n740), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U795 ( .A1(n752), .A2(G469), .ZN(n746) );
  XOR2_X1 U796 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n743) );
  XNOR2_X1 U797 ( .A(n743), .B(KEYINPUT122), .ZN(n744) );
  XNOR2_X1 U798 ( .A(n742), .B(n744), .ZN(n745) );
  XNOR2_X1 U799 ( .A(n746), .B(n745), .ZN(n747) );
  NOR2_X1 U800 ( .A1(n757), .A2(n747), .ZN(G54) );
  NAND2_X1 U801 ( .A1(n752), .A2(G478), .ZN(n750) );
  XOR2_X1 U802 ( .A(KEYINPUT124), .B(n748), .Z(n749) );
  XNOR2_X1 U803 ( .A(n750), .B(n749), .ZN(n751) );
  NOR2_X1 U804 ( .A1(n757), .A2(n751), .ZN(G63) );
  NAND2_X1 U805 ( .A1(n752), .A2(G217), .ZN(n755) );
  XNOR2_X1 U806 ( .A(n753), .B(KEYINPUT125), .ZN(n754) );
  XNOR2_X1 U807 ( .A(n755), .B(n754), .ZN(n756) );
  NOR2_X1 U808 ( .A1(n757), .A2(n756), .ZN(G66) );
  NAND2_X1 U809 ( .A1(G953), .A2(G224), .ZN(n758) );
  XNOR2_X1 U810 ( .A(KEYINPUT61), .B(n758), .ZN(n759) );
  NAND2_X1 U811 ( .A1(n759), .A2(G898), .ZN(n760) );
  NAND2_X1 U812 ( .A1(n761), .A2(n760), .ZN(n767) );
  XOR2_X1 U813 ( .A(G101), .B(KEYINPUT126), .Z(n762) );
  XNOR2_X1 U814 ( .A(n763), .B(n762), .ZN(n765) );
  NAND2_X1 U815 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U816 ( .A(n767), .B(n766), .Z(G69) );
  XNOR2_X1 U817 ( .A(n768), .B(KEYINPUT127), .ZN(n770) );
  XNOR2_X1 U818 ( .A(n770), .B(n769), .ZN(n771) );
  XOR2_X1 U819 ( .A(n772), .B(n771), .Z(n776) );
  XNOR2_X1 U820 ( .A(n773), .B(n776), .ZN(n775) );
  NAND2_X1 U821 ( .A1(n775), .A2(n774), .ZN(n780) );
  XNOR2_X1 U822 ( .A(G227), .B(n776), .ZN(n777) );
  NAND2_X1 U823 ( .A1(n777), .A2(G900), .ZN(n778) );
  NAND2_X1 U824 ( .A1(n778), .A2(G953), .ZN(n779) );
  NAND2_X1 U825 ( .A1(n780), .A2(n779), .ZN(G72) );
  XNOR2_X1 U826 ( .A(G119), .B(n781), .ZN(G21) );
  XNOR2_X1 U827 ( .A(n782), .B(KEYINPUT118), .ZN(n783) );
  XNOR2_X1 U828 ( .A(n783), .B(KEYINPUT37), .ZN(n784) );
  XNOR2_X1 U829 ( .A(G125), .B(n784), .ZN(G27) );
  XNOR2_X1 U830 ( .A(G131), .B(n785), .ZN(G33) );
  XNOR2_X1 U831 ( .A(G137), .B(n786), .ZN(G39) );
endmodule

