//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(G134), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G137), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n187), .A2(G137), .ZN(new_n190));
  OAI21_X1  g004(.A(G131), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT11), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n192), .B1(new_n187), .B2(G137), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n194), .A2(KEYINPUT11), .A3(G134), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n193), .A2(new_n195), .A3(new_n196), .A4(new_n188), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n202), .A2(KEYINPUT1), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  AND3_X1   g018(.A1(new_n204), .A2(KEYINPUT66), .A3(G146), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT66), .B1(new_n204), .B2(G146), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n201), .B(new_n203), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT69), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT1), .ZN(new_n209));
  AOI21_X1  g023(.A(new_n209), .B1(G143), .B2(new_n200), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n204), .A2(G146), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n200), .A2(G143), .ZN(new_n212));
  OAI22_X1  g026(.A1(new_n210), .A2(new_n202), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n207), .A2(new_n208), .A3(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n208), .B1(new_n207), .B2(new_n213), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n199), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT2), .B(G113), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(KEYINPUT67), .A2(G119), .ZN(new_n219));
  INV_X1    g033(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(KEYINPUT67), .A2(G119), .ZN(new_n221));
  OAI21_X1  g035(.A(G116), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G119), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n223), .A2(G116), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n218), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G116), .ZN(new_n228));
  OR2_X1    g042(.A1(KEYINPUT67), .A2(G119), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(new_n219), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT68), .B1(new_n230), .B2(new_n224), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n222), .A2(new_n232), .A3(new_n225), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n227), .B1(new_n234), .B2(new_n217), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n193), .A2(new_n188), .A3(new_n195), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G131), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(new_n197), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n204), .A2(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n201), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT64), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT0), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n242), .A2(new_n243), .A3(new_n202), .ZN(new_n244));
  OAI21_X1  g058(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n240), .A2(new_n241), .A3(new_n244), .A4(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT65), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT66), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n248), .B1(new_n200), .B2(G143), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n204), .A2(KEYINPUT66), .A3(G146), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n211), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT0), .A3(G128), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n245), .A2(new_n241), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT65), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n253), .A2(new_n254), .A3(new_n244), .A4(new_n240), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n238), .A2(new_n247), .A3(new_n252), .A4(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n216), .A2(new_n235), .A3(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n235), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n207), .A2(new_n213), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n199), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n216), .A2(new_n235), .A3(KEYINPUT28), .A4(new_n256), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n259), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(G237), .A2(G953), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G210), .ZN(new_n268));
  XNOR2_X1  g082(.A(new_n268), .B(G101), .ZN(new_n269));
  XNOR2_X1  g083(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT70), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n266), .A2(new_n275), .A3(new_n272), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT30), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n263), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n216), .A2(KEYINPUT30), .A3(new_n256), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n278), .A2(new_n279), .A3(new_n260), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n257), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT31), .B1(new_n281), .B2(new_n272), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT31), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n280), .A2(new_n283), .A3(new_n257), .A4(new_n271), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n274), .A2(new_n276), .A3(new_n282), .A4(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(G472), .A2(G902), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n285), .A2(KEYINPUT32), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT72), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n261), .A2(KEYINPUT69), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n207), .A2(new_n213), .A3(new_n208), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n198), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n256), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n260), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  AND2_X1   g107(.A1(new_n271), .A2(KEYINPUT29), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n259), .A2(new_n265), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(KEYINPUT29), .B1(new_n281), .B2(new_n272), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n259), .A2(new_n264), .A3(new_n265), .A4(new_n271), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G472), .ZN(new_n301));
  OAI21_X1  g115(.A(KEYINPUT71), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT71), .ZN(new_n303));
  INV_X1    g117(.A(new_n299), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n271), .B1(new_n280), .B2(new_n257), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n304), .A2(new_n305), .A3(KEYINPUT29), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n303), .B(G472), .C1(new_n306), .C2(new_n297), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n285), .A2(new_n286), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT32), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT72), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n285), .A2(new_n312), .A3(KEYINPUT32), .A4(new_n286), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n288), .A2(new_n308), .A3(new_n311), .A4(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT77), .ZN(new_n315));
  INV_X1    g129(.A(G953), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n316), .A2(G221), .A3(G234), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(G137), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT73), .B(KEYINPUT22), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n322), .A2(KEYINPUT16), .A3(G140), .ZN(new_n323));
  XNOR2_X1  g137(.A(G125), .B(G140), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(KEYINPUT16), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n325), .B(G146), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT23), .ZN(new_n327));
  XNOR2_X1  g141(.A(KEYINPUT67), .B(G119), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n327), .B1(new_n328), .B2(G128), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n223), .A2(G128), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n330), .B1(new_n328), .B2(G128), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n329), .B1(new_n331), .B2(new_n327), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G110), .ZN(new_n333));
  XOR2_X1   g147(.A(KEYINPUT24), .B(G110), .Z(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  AND3_X1   g149(.A1(new_n326), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n325), .A2(G146), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n324), .A2(new_n200), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(G110), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n340), .B(new_n329), .C1(new_n331), .C2(new_n327), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n331), .A2(new_n334), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n339), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n321), .B1(new_n336), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n344), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n326), .A2(new_n333), .A3(new_n335), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(new_n320), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G217), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n350), .B1(G234), .B2(new_n296), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n351), .A2(G902), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(KEYINPUT75), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n349), .A2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT76), .ZN(new_n356));
  NOR3_X1   g170(.A1(new_n336), .A2(new_n344), .A3(new_n321), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n320), .B1(new_n346), .B2(new_n347), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n296), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT74), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT25), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(KEYINPUT25), .ZN(new_n362));
  OR2_X1    g176(.A1(new_n360), .A2(KEYINPUT25), .ZN(new_n363));
  NAND4_X1  g177(.A1(new_n349), .A2(new_n296), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n351), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n356), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n314), .A2(new_n315), .A3(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n315), .B1(new_n314), .B2(new_n367), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(G237), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(new_n316), .A3(G214), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT85), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(G143), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n267), .B(G214), .C1(new_n373), .C2(G143), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(KEYINPUT18), .A2(G131), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(KEYINPUT86), .B1(new_n324), .B2(new_n200), .ZN(new_n380));
  OR3_X1    g194(.A1(new_n380), .A2(new_n200), .A3(new_n324), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n380), .B1(new_n200), .B2(new_n324), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n379), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT87), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n324), .A2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n385), .B(KEYINPUT19), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(G146), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n377), .A2(G131), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n375), .A2(new_n376), .A3(new_n196), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n337), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n383), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  XNOR2_X1  g206(.A(G113), .B(G122), .ZN(new_n393));
  INV_X1    g207(.A(G104), .ZN(new_n394));
  XNOR2_X1  g208(.A(new_n393), .B(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT17), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n388), .A2(new_n398), .A3(new_n389), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT88), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n325), .B(new_n200), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n377), .A2(KEYINPUT17), .A3(G131), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT88), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n388), .A2(new_n403), .A3(new_n398), .A4(new_n389), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n400), .A2(new_n401), .A3(new_n402), .A4(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(new_n383), .A3(new_n395), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n397), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G475), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(new_n408), .A3(new_n296), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n409), .B(KEYINPUT20), .Z(new_n410));
  INV_X1    g224(.A(KEYINPUT89), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n405), .A2(new_n383), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n411), .B1(new_n412), .B2(new_n396), .ZN(new_n413));
  AOI211_X1 g227(.A(KEYINPUT89), .B(new_n395), .C1(new_n405), .C2(new_n383), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n406), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT90), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n415), .A2(new_n416), .A3(new_n296), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n416), .B1(new_n415), .B2(new_n296), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n410), .B1(new_n419), .B2(G475), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT94), .ZN(new_n421));
  NAND2_X1  g235(.A1(G234), .A2(G237), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n422), .A2(G952), .A3(new_n316), .ZN(new_n423));
  XOR2_X1   g237(.A(KEYINPUT21), .B(G898), .Z(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n422), .A2(G902), .A3(G953), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n423), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(G116), .B(G122), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT14), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n228), .A2(KEYINPUT14), .A3(G122), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(G107), .A3(new_n432), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n433), .A2(KEYINPUT92), .ZN(new_n434));
  INV_X1    g248(.A(G107), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n433), .B2(KEYINPUT92), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT91), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n438), .B1(new_n204), .B2(G128), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n202), .A2(KEYINPUT91), .A3(G143), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n439), .A2(new_n440), .B1(G128), .B2(new_n204), .ZN(new_n441));
  OR2_X1    g255(.A1(new_n441), .A2(G134), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(G134), .ZN(new_n443));
  NAND4_X1  g257(.A1(new_n434), .A2(new_n437), .A3(new_n442), .A4(new_n443), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT13), .B1(new_n439), .B2(new_n440), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n445), .A2(new_n187), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n446), .A2(new_n441), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n441), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n429), .A2(new_n435), .ZN(new_n449));
  OAI22_X1  g263(.A1(new_n447), .A2(new_n448), .B1(new_n449), .B2(new_n436), .ZN(new_n450));
  XOR2_X1   g264(.A(KEYINPUT9), .B(G234), .Z(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NOR3_X1   g266(.A1(new_n452), .A2(new_n350), .A3(G953), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n444), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n453), .B1(new_n444), .B2(new_n450), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n296), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT15), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n456), .A2(new_n457), .A3(G478), .ZN(new_n458));
  INV_X1    g272(.A(G478), .ZN(new_n459));
  OAI221_X1 g273(.A(new_n296), .B1(KEYINPUT15), .B2(new_n459), .C1(new_n454), .C2(new_n455), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n458), .A2(KEYINPUT93), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT93), .B1(new_n458), .B2(new_n460), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n420), .A2(new_n421), .A3(new_n428), .A4(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n415), .A2(new_n296), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT90), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n415), .A2(new_n416), .A3(new_n296), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(G475), .A3(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n409), .B(KEYINPUT20), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n428), .A4(new_n463), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(KEYINPUT94), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(KEYINPUT3), .B1(new_n394), .B2(G107), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT3), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n474), .A2(new_n435), .A3(G104), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n394), .A2(G107), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(KEYINPUT79), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT79), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n473), .A2(new_n475), .A3(new_n479), .A4(new_n476), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n478), .A2(G101), .A3(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G101), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n473), .A2(new_n475), .A3(new_n482), .A4(new_n476), .ZN(new_n483));
  AND2_X1   g297(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT4), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n478), .A2(new_n486), .A3(G101), .A4(new_n480), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n218), .B1(new_n231), .B2(new_n233), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n485), .B(new_n487), .C1(new_n488), .C2(new_n227), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n231), .A2(KEYINPUT5), .A3(new_n233), .ZN(new_n490));
  INV_X1    g304(.A(G113), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT5), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n491), .B1(new_n230), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n476), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n394), .A2(G107), .ZN(new_n496));
  OAI21_X1  g310(.A(G101), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n483), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n494), .A2(new_n226), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n489), .A2(new_n500), .ZN(new_n501));
  XOR2_X1   g315(.A(G110), .B(G122), .Z(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n502), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n489), .A2(new_n500), .A3(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n503), .A2(KEYINPUT6), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT6), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n501), .A2(new_n507), .A3(new_n502), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n261), .A2(G125), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n247), .A2(new_n252), .A3(new_n255), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(G125), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n316), .A2(G224), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n506), .A2(new_n508), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n510), .A2(G125), .ZN(new_n515));
  INV_X1    g329(.A(new_n509), .ZN(new_n516));
  NAND2_X1  g330(.A1(KEYINPUT83), .A2(KEYINPUT7), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n515), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n512), .A2(KEYINPUT7), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n511), .A2(new_n517), .A3(new_n519), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n222), .A2(KEYINPUT5), .A3(new_n225), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n493), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n498), .B1(new_n524), .B2(new_n226), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n227), .B1(new_n490), .B2(new_n493), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n525), .B1(new_n526), .B2(new_n498), .ZN(new_n527));
  XOR2_X1   g341(.A(KEYINPUT82), .B(KEYINPUT8), .Z(new_n528));
  XNOR2_X1  g342(.A(new_n502), .B(new_n528), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n521), .A2(new_n522), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(G902), .B1(new_n530), .B2(new_n505), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n514), .A2(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(G210), .B1(G237), .B2(G902), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n514), .A2(new_n531), .A3(new_n533), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(KEYINPUT84), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT84), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n532), .A2(new_n538), .A3(new_n534), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(G214), .B1(G237), .B2(G902), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n201), .B1(new_n205), .B2(new_n206), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n202), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT80), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n544), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT80), .B1(new_n251), .B2(new_n545), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n549), .A3(new_n207), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n499), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT10), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n510), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(new_n485), .A3(new_n487), .ZN(new_n555));
  OAI211_X1 g369(.A(KEYINPUT10), .B(new_n499), .C1(new_n214), .C2(new_n215), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n238), .ZN(new_n558));
  INV_X1    g372(.A(new_n238), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n553), .A2(new_n555), .A3(new_n559), .A4(new_n556), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n316), .A2(G227), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(G140), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT78), .B(G110), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n498), .A2(new_n213), .A3(new_n207), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n559), .B1(new_n551), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g382(.A(KEYINPUT81), .B1(new_n568), .B2(KEYINPUT12), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT81), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT12), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n499), .A2(new_n261), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n572), .B1(new_n499), .B2(new_n550), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n570), .B(new_n571), .C1(new_n573), .C2(new_n559), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n568), .A2(KEYINPUT12), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n569), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n565), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n560), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n566), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G469), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n581), .A3(new_n296), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n576), .A2(new_n560), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n565), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n578), .A2(new_n558), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(G469), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(G469), .A2(G902), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(G221), .B1(new_n452), .B2(G902), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n472), .A2(new_n543), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n370), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(new_n482), .ZN(G3));
  INV_X1    g407(.A(KEYINPUT99), .ZN(new_n594));
  AND2_X1   g408(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n595));
  NOR2_X1   g409(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n454), .A2(new_n455), .A3(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n444), .A2(new_n450), .ZN(new_n599));
  INV_X1    g413(.A(new_n453), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n444), .A2(new_n450), .A3(new_n453), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n595), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(G478), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  OR2_X1    g418(.A1(new_n456), .A2(G478), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n459), .A2(new_n296), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n604), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(KEYINPUT98), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT98), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n604), .A2(new_n605), .A3(new_n610), .A4(new_n607), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n417), .A2(new_n418), .A3(new_n408), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n612), .B1(new_n613), .B2(new_n410), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT96), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n535), .A2(new_n615), .A3(new_n536), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n533), .B1(new_n514), .B2(new_n531), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n542), .B1(new_n617), .B2(KEYINPUT96), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n428), .A3(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n594), .B1(new_n614), .B2(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n616), .A2(new_n428), .A3(new_n618), .ZN(new_n621));
  AOI22_X1  g435(.A1(new_n468), .A2(new_n469), .B1(new_n609), .B2(new_n611), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(KEYINPUT99), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n301), .B1(new_n285), .B2(new_n296), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT95), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(KEYINPUT95), .B1(new_n285), .B2(new_n286), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n627), .B1(new_n625), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n588), .A2(new_n589), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n629), .A2(new_n366), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT34), .B(G104), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  NAND2_X1  g448(.A1(new_n468), .A2(new_n469), .ZN(new_n635));
  NOR3_X1   g449(.A1(new_n619), .A2(new_n635), .A3(new_n463), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(KEYINPUT35), .B(G107), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(G9));
  NAND2_X1  g453(.A1(new_n346), .A2(new_n347), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n320), .A2(KEYINPUT36), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(new_n354), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n365), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(KEYINPUT100), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n629), .A2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n472), .A2(new_n543), .A3(new_n590), .A4(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT37), .B(G110), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT101), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n647), .B(new_n649), .ZN(G12));
  NAND2_X1  g464(.A1(new_n616), .A2(new_n618), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n644), .B(new_n653), .ZN(new_n654));
  AND4_X1   g468(.A1(new_n314), .A2(new_n590), .A3(new_n652), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(KEYINPUT102), .B(G900), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n423), .B1(new_n426), .B2(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n635), .A2(new_n463), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G128), .ZN(G30));
  INV_X1    g474(.A(KEYINPUT38), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n540), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n537), .A2(KEYINPUT38), .A3(new_n539), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n281), .A2(new_n271), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n293), .A2(new_n257), .A3(new_n272), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n665), .A2(new_n296), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n667), .A2(G472), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n288), .A2(new_n311), .A3(new_n313), .A4(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n420), .A2(new_n463), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n664), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n657), .B(KEYINPUT39), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n590), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n671), .B1(new_n675), .B2(KEYINPUT40), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n644), .A2(new_n542), .ZN(new_n677));
  OAI211_X1 g491(.A(new_n676), .B(new_n677), .C1(KEYINPUT40), .C2(new_n675), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  INV_X1    g493(.A(new_n657), .ZN(new_n680));
  AND3_X1   g494(.A1(new_n635), .A2(new_n612), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n655), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  NAND2_X1  g497(.A1(new_n580), .A2(new_n296), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G469), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n589), .A3(new_n582), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  AND3_X1   g501(.A1(new_n314), .A2(new_n367), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n624), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND2_X1  g505(.A1(new_n688), .A2(new_n636), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  NOR3_X1   g507(.A1(new_n645), .A2(new_n651), .A3(new_n686), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n472), .A2(new_n314), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G119), .ZN(G21));
  NAND3_X1  g510(.A1(new_n259), .A2(new_n265), .A3(new_n293), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n697), .A2(new_n272), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n282), .A2(new_n284), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n625), .B1(new_n286), .B2(new_n699), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n700), .A2(new_n367), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n701), .A2(new_n621), .A3(new_n670), .A4(new_n687), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G122), .ZN(G24));
  AND2_X1   g517(.A1(new_n700), .A2(new_n644), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n686), .A2(new_n651), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n704), .A2(new_n622), .A3(new_n680), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G125), .ZN(G27));
  INV_X1    g521(.A(KEYINPUT106), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n588), .A2(KEYINPUT104), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n582), .A2(new_n586), .A3(new_n710), .A4(new_n587), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n709), .A2(new_n589), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n536), .A2(KEYINPUT84), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n617), .ZN(new_n714));
  INV_X1    g528(.A(new_n539), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n541), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT105), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n540), .A2(new_n718), .A3(new_n541), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n712), .A2(new_n717), .A3(new_n681), .A4(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n314), .A2(new_n367), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n708), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n718), .B1(new_n540), .B2(new_n541), .ZN(new_n723));
  AOI211_X1 g537(.A(KEYINPUT105), .B(new_n542), .C1(new_n537), .C2(new_n539), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n635), .A2(new_n612), .A3(new_n680), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n721), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(KEYINPUT106), .A3(new_n727), .A4(new_n712), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT42), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n722), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n308), .A2(new_n287), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n366), .B1(new_n731), .B2(new_n311), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n726), .A2(KEYINPUT42), .A3(new_n712), .A4(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G131), .ZN(G33));
  NOR2_X1   g549(.A1(new_n723), .A2(new_n724), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n727), .A2(new_n736), .A3(new_n658), .A4(new_n712), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT107), .B(G134), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(G36));
  NAND2_X1  g553(.A1(new_n584), .A2(new_n585), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT45), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(G469), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT108), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n584), .A2(KEYINPUT45), .A3(new_n585), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT108), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n742), .A2(new_n746), .A3(G469), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n744), .A2(new_n745), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n587), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT109), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n749), .A2(new_n750), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n748), .A2(new_n753), .A3(KEYINPUT46), .A4(new_n587), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n751), .A2(new_n752), .A3(new_n582), .A4(new_n754), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(new_n589), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n672), .A3(new_n736), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n420), .A2(new_n612), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT43), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT43), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n420), .A2(new_n760), .A3(new_n612), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n759), .A2(new_n629), .A3(new_n644), .A4(new_n761), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT44), .Z(new_n763));
  OR2_X1    g577(.A1(new_n757), .A2(new_n763), .ZN(new_n764));
  XOR2_X1   g578(.A(KEYINPUT110), .B(G137), .Z(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G39));
  NAND2_X1  g580(.A1(new_n755), .A2(new_n589), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT47), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n755), .A2(KEYINPUT47), .A3(new_n589), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n314), .A2(new_n367), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n771), .A2(new_n726), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(G140), .ZN(G42));
  INV_X1    g588(.A(new_n589), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n366), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n685), .A2(new_n582), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT111), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT49), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n780), .A2(new_n542), .A3(new_n758), .ZN(new_n781));
  XOR2_X1   g595(.A(new_n781), .B(KEYINPUT112), .Z(new_n782));
  AOI21_X1  g596(.A(new_n669), .B1(new_n778), .B2(new_n779), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n782), .A2(new_n663), .A3(new_n662), .A4(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n778), .A2(new_n775), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n769), .A2(new_n770), .A3(new_n786), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n759), .A2(new_n701), .A3(new_n423), .A4(new_n761), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(new_n736), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT115), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n759), .A2(new_n423), .A3(new_n761), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n662), .A2(new_n663), .A3(new_n687), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n793), .A2(new_n542), .A3(new_n795), .A4(new_n701), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT50), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n792), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n788), .A2(new_n541), .A3(new_n794), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n799), .A2(new_n801), .A3(KEYINPUT50), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT114), .B1(new_n796), .B2(new_n797), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n798), .B(new_n800), .C1(new_n802), .C2(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n723), .A2(new_n724), .A3(new_n686), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n793), .A2(new_n704), .A3(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n669), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n805), .A2(new_n367), .A3(new_n423), .A4(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n420), .A2(new_n609), .A3(new_n611), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n804), .A2(new_n806), .A3(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n785), .B1(new_n791), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT117), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n798), .A2(new_n800), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n801), .B1(new_n799), .B2(KEYINPUT50), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n796), .A2(KEYINPUT114), .A3(new_n797), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n810), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n816), .B1(new_n821), .B2(new_n806), .ZN(new_n822));
  AND4_X1   g636(.A1(new_n816), .A2(new_n804), .A3(new_n806), .A4(new_n811), .ZN(new_n823));
  OAI211_X1 g637(.A(KEYINPUT51), .B(new_n790), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(KEYINPUT116), .B(new_n785), .C1(new_n791), .C2(new_n812), .ZN(new_n825));
  OAI211_X1 g639(.A(G952), .B(new_n316), .C1(new_n808), .C2(new_n614), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n793), .A2(new_n732), .A3(new_n805), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n827), .A2(KEYINPUT48), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(KEYINPUT48), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n815), .A2(new_n824), .A3(new_n825), .A4(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n788), .A2(new_n651), .A3(new_n686), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n458), .A2(new_n460), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n314), .A2(new_n590), .A3(new_n654), .A4(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n622), .A2(new_n700), .A3(new_n644), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n709), .A2(new_n589), .A3(new_n711), .ZN(new_n837));
  OAI22_X1  g651(.A1(new_n835), .A2(new_n635), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n838), .A2(new_n680), .A3(new_n736), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n614), .B1(new_n834), .B2(new_n635), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n631), .A2(new_n543), .A3(new_n428), .A4(new_n840), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n647), .B(new_n841), .C1(new_n370), .C2(new_n591), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n689), .A2(new_n695), .A3(new_n692), .A4(new_n702), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n839), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n737), .B1(new_n730), .B2(new_n733), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n655), .B1(new_n658), .B2(new_n681), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n420), .A2(new_n651), .A3(new_n463), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n644), .A2(new_n657), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n712), .A2(new_n847), .A3(new_n669), .A4(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n846), .A2(new_n706), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT113), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n850), .A2(new_n851), .A3(KEYINPUT52), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n844), .A2(new_n845), .A3(new_n854), .A4(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n850), .B(new_n853), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(KEYINPUT53), .A3(new_n844), .A4(new_n845), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n833), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n856), .A2(KEYINPUT53), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n859), .A2(new_n857), .A3(new_n844), .A4(new_n845), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT54), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n831), .A2(new_n832), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(G952), .A2(G953), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n784), .B1(new_n866), .B2(new_n867), .ZN(G75));
  OR2_X1    g682(.A1(new_n316), .A2(G952), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT118), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n862), .A2(G210), .A3(G902), .A4(new_n863), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT56), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n506), .A2(new_n508), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n873), .B(new_n513), .Z(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(KEYINPUT55), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n871), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n875), .B1(new_n871), .B2(new_n872), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n870), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n878), .B(new_n879), .ZN(G51));
  INV_X1    g694(.A(new_n870), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n862), .A2(KEYINPUT54), .A3(new_n863), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT121), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n862), .A2(new_n863), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n833), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n862), .A2(new_n886), .A3(KEYINPUT54), .A4(new_n863), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n883), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n587), .B(KEYINPUT120), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n889), .B(KEYINPUT57), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n580), .B(KEYINPUT122), .Z(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OR3_X1    g707(.A1(new_n884), .A2(new_n296), .A3(new_n748), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n881), .B1(new_n893), .B2(new_n894), .ZN(G54));
  AND2_X1   g709(.A1(new_n862), .A2(new_n863), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(new_n407), .Z(new_n898));
  NOR2_X1   g712(.A1(new_n898), .A2(new_n881), .ZN(G60));
  XNOR2_X1  g713(.A(KEYINPUT124), .B(KEYINPUT59), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n607), .B(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n901), .B1(new_n861), .B2(new_n864), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n598), .A2(new_n603), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT123), .Z(new_n904));
  AOI21_X1  g718(.A(new_n881), .B1(new_n902), .B2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n901), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n888), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT125), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n905), .A2(new_n908), .A3(KEYINPUT125), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(G63));
  INV_X1    g727(.A(KEYINPUT60), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n350), .B2(new_n296), .ZN(new_n915));
  NAND3_X1  g729(.A1(KEYINPUT60), .A2(G217), .A3(G902), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n896), .A2(new_n642), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n884), .B1(new_n915), .B2(new_n916), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n918), .B(new_n870), .C1(new_n919), .C2(new_n349), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT61), .Z(G66));
  INV_X1    g735(.A(G224), .ZN(new_n922));
  OAI21_X1  g736(.A(G953), .B1(new_n425), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n842), .A2(new_n843), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n923), .B1(new_n924), .B2(G953), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n873), .B1(G898), .B2(new_n316), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n925), .B(new_n926), .ZN(G69));
  AND2_X1   g741(.A1(new_n846), .A2(new_n706), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n928), .B1(new_n757), .B2(new_n763), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(KEYINPUT127), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT127), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n931), .B(new_n928), .C1(new_n757), .C2(new_n763), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n756), .A2(new_n672), .A3(new_n732), .A4(new_n847), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n934), .A2(new_n845), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n933), .A2(new_n935), .A3(new_n316), .A4(new_n773), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n278), .A2(new_n279), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n937), .B(new_n386), .ZN(new_n938));
  NAND2_X1  g752(.A1(G900), .A2(G953), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n938), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n678), .A2(new_n928), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT62), .B1(new_n678), .B2(new_n928), .ZN(new_n945));
  INV_X1    g759(.A(new_n370), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n736), .A3(new_n840), .ZN(new_n947));
  OAI22_X1  g761(.A1(new_n944), .A2(new_n945), .B1(new_n675), .B2(new_n947), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n764), .A2(new_n773), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n941), .B1(new_n950), .B2(G953), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n940), .A2(KEYINPUT126), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n316), .B1(G227), .B2(G900), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n953), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n940), .A2(KEYINPUT126), .A3(new_n955), .A4(new_n951), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(G72));
  NAND2_X1  g771(.A1(new_n950), .A2(new_n924), .ZN(new_n958));
  NAND2_X1  g772(.A1(G472), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT63), .Z(new_n960));
  AOI21_X1  g774(.A(new_n665), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n280), .A2(new_n257), .A3(new_n272), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n933), .A2(new_n935), .A3(new_n773), .A4(new_n924), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n963), .B2(new_n960), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n858), .A2(new_n860), .ZN(new_n965));
  AND4_X1   g779(.A1(new_n665), .A2(new_n965), .A3(new_n960), .A4(new_n962), .ZN(new_n966));
  NOR4_X1   g780(.A1(new_n961), .A2(new_n964), .A3(new_n881), .A4(new_n966), .ZN(G57));
endmodule


