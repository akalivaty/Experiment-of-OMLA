//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n561, new_n562, new_n563, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1232, new_n1233;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(new_n459), .A2(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(new_n459), .ZN(new_n463));
  INV_X1    g038(.A(G137), .ZN(new_n464));
  OAI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(G125), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n459), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n465), .A2(new_n468), .ZN(G160));
  OR2_X1    g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n459), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G124), .ZN(new_n473));
  OR2_X1    g048(.A1(G100), .A2(G2105), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n474), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n475));
  INV_X1    g050(.A(G136), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n473), .B(new_n475), .C1(new_n476), .C2(new_n463), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G162));
  INV_X1    g053(.A(G138), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G2105), .ZN(new_n480));
  AND2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  NOR2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(KEYINPUT4), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n480), .B(new_n485), .C1(new_n482), .C2(new_n481), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n488));
  OR2_X1    g063(.A1(new_n459), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n472), .A2(G126), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n487), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n488), .B1(new_n487), .B2(new_n492), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n493), .A2(new_n494), .ZN(G164));
  AND2_X1   g070(.A1(KEYINPUT6), .A2(G651), .ZN(new_n496));
  NOR2_X1   g071(.A1(KEYINPUT6), .A2(G651), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  AND2_X1   g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NOR2_X1   g074(.A1(KEYINPUT5), .A2(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g076(.A(KEYINPUT67), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT5), .B(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n503), .B(new_n504), .C1(new_n497), .C2(new_n496), .ZN(new_n505));
  AND3_X1   g080(.A1(new_n502), .A2(new_n505), .A3(G88), .ZN(new_n506));
  INV_X1    g081(.A(G75), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  OAI21_X1  g083(.A(KEYINPUT68), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(G75), .A3(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G62), .ZN(new_n513));
  OR2_X1    g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OAI21_X1  g091(.A(G651), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n498), .A2(new_n508), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(KEYINPUT69), .B1(new_n506), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n509), .B(new_n511), .C1(new_n501), .C2(new_n513), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n522), .A2(G651), .B1(new_n518), .B2(G50), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT69), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n502), .A2(new_n505), .ZN(new_n526));
  OAI211_X1 g101(.A(new_n523), .B(new_n524), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n521), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n518), .A2(G51), .B1(new_n503), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n502), .A2(new_n505), .A3(G89), .ZN(new_n532));
  NAND3_X1  g107(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n533));
  XNOR2_X1  g108(.A(new_n533), .B(KEYINPUT7), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT70), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(KEYINPUT70), .B1(new_n532), .B2(new_n534), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n531), .B1(new_n537), .B2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  AND2_X1   g115(.A1(new_n502), .A2(new_n505), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G90), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  INV_X1    g118(.A(G77), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n501), .A2(new_n543), .B1(new_n544), .B2(new_n508), .ZN(new_n545));
  INV_X1    g120(.A(KEYINPUT71), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  OAI221_X1 g122(.A(KEYINPUT71), .B1(new_n544), .B2(new_n508), .C1(new_n501), .C2(new_n543), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n547), .A2(G651), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n518), .A2(G52), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n542), .A2(new_n549), .A3(new_n550), .ZN(G171));
  NAND2_X1  g126(.A1(new_n541), .A2(G81), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n501), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n555), .A2(G651), .B1(new_n518), .B2(G43), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(new_n557));
  INV_X1    g132(.A(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G860), .ZN(G153));
  NAND4_X1  g134(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g135(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n561));
  NAND2_X1  g136(.A1(G1), .A2(G3), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n561), .B(new_n562), .ZN(new_n563));
  NAND4_X1  g138(.A1(G319), .A2(G483), .A3(G661), .A4(new_n563), .ZN(G188));
  OAI211_X1 g139(.A(G53), .B(G543), .C1(new_n496), .C2(new_n497), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT9), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n566), .A2(KEYINPUT73), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n565), .B(new_n567), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n502), .A2(new_n505), .A3(G91), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n501), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n568), .A2(new_n569), .A3(new_n573), .ZN(G299));
  NAND3_X1  g149(.A1(new_n542), .A2(new_n549), .A3(new_n550), .ZN(G301));
  NAND2_X1  g150(.A1(new_n541), .A2(G87), .ZN(new_n576));
  OR2_X1    g151(.A1(new_n503), .A2(G74), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n577), .A2(G651), .B1(new_n518), .B2(G49), .ZN(new_n578));
  AND2_X1   g153(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G288));
  NAND2_X1  g155(.A1(new_n541), .A2(G86), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n501), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n584), .A2(G651), .B1(new_n518), .B2(G48), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n581), .A2(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(G72), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G60), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n501), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n589), .A2(G651), .B1(new_n518), .B2(G47), .ZN(new_n590));
  INV_X1    g165(.A(G85), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n526), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n593));
  XNOR2_X1  g168(.A(new_n592), .B(new_n593), .ZN(G290));
  INV_X1    g169(.A(G868), .ZN(new_n595));
  OR3_X1    g170(.A1(G171), .A2(KEYINPUT75), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(KEYINPUT75), .B1(G171), .B2(new_n595), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT76), .ZN(new_n599));
  XNOR2_X1  g174(.A(KEYINPUT77), .B(G66), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n501), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n518), .A2(G54), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n541), .A2(KEYINPUT10), .A3(G92), .ZN(new_n605));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n526), .B2(new_n607), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n604), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  OAI211_X1 g184(.A(new_n596), .B(new_n597), .C1(G868), .C2(new_n609), .ZN(G284));
  OAI211_X1 g185(.A(new_n596), .B(new_n597), .C1(G868), .C2(new_n609), .ZN(G321));
  NAND2_X1  g186(.A1(G299), .A2(new_n595), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G168), .B2(new_n595), .ZN(G297));
  OAI21_X1  g188(.A(new_n612), .B1(G168), .B2(new_n595), .ZN(G280));
  XNOR2_X1  g189(.A(KEYINPUT78), .B(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n609), .B1(G860), .B2(new_n615), .ZN(G148));
  NAND2_X1  g191(.A1(new_n609), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(G868), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n618), .B1(G868), .B2(new_n558), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n462), .A2(new_n460), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XOR2_X1   g198(.A(KEYINPUT79), .B(G2100), .Z(new_n624));
  OR2_X1    g199(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n624), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n472), .A2(G123), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n459), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  INV_X1    g204(.A(G135), .ZN(new_n630));
  OAI221_X1 g205(.A(new_n627), .B1(new_n628), .B2(new_n629), .C1(new_n630), .C2(new_n463), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(G2096), .Z(new_n632));
  NAND3_X1  g207(.A1(new_n625), .A2(new_n626), .A3(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT80), .ZN(G156));
  XOR2_X1   g209(.A(G2451), .B(G2454), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT16), .ZN(new_n636));
  XNOR2_X1  g211(.A(G1341), .B(G1348), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT81), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n643), .B2(new_n642), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n639), .B(new_n645), .Z(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(G14), .A3(new_n649), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(G401));
  XNOR2_X1  g226(.A(G2084), .B(G2090), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT82), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G2067), .B(G2678), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT83), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2072), .B(G2078), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT17), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n654), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n656), .B2(new_n657), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT84), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NAND3_X1  g237(.A1(new_n654), .A2(new_n656), .A3(new_n657), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT18), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n656), .A2(new_n653), .A3(new_n658), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2096), .B(G2100), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G227));
  XOR2_X1   g245(.A(G1991), .B(G1996), .Z(new_n671));
  XNOR2_X1  g246(.A(G1971), .B(G1976), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT19), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  NOR2_X1   g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n675), .A2(new_n676), .ZN(new_n679));
  NOR3_X1   g254(.A1(new_n674), .A2(new_n679), .A3(new_n677), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n674), .A2(new_n679), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT85), .B(KEYINPUT20), .Z(new_n682));
  AOI211_X1 g257(.A(new_n678), .B(new_n680), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n684));
  OR2_X1    g259(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n684), .B1(new_n683), .B2(new_n685), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n671), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n688), .ZN(new_n690));
  INV_X1    g265(.A(new_n671), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n690), .A2(new_n686), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n694), .B(KEYINPUT87), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XOR2_X1   g271(.A(new_n695), .B(new_n696), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n693), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n689), .A2(new_n692), .A3(new_n697), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(G229));
  NAND2_X1  g276(.A1(G168), .A2(G16), .ZN(new_n702));
  OR2_X1    g277(.A1(G16), .A2(G21), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT100), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(G1966), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT30), .B(G28), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  OR2_X1    g283(.A1(KEYINPUT31), .A2(G11), .ZN(new_n709));
  NAND2_X1  g284(.A1(KEYINPUT31), .A2(G11), .ZN(new_n710));
  AOI22_X1  g285(.A1(new_n707), .A2(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n711), .B1(new_n631), .B2(new_n708), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT24), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n708), .B1(new_n713), .B2(G34), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n713), .B2(G34), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(G160), .B2(G29), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n712), .B1(new_n716), .B2(G2084), .ZN(new_n717));
  INV_X1    g292(.A(G16), .ZN(new_n718));
  NOR2_X1   g293(.A1(G171), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G5), .B2(new_n718), .ZN(new_n720));
  INV_X1    g295(.A(G1961), .ZN(new_n721));
  OAI221_X1 g296(.A(new_n717), .B1(G2084), .B2(new_n716), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n708), .A2(G32), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n472), .A2(G129), .ZN(new_n724));
  XOR2_X1   g299(.A(new_n724), .B(KEYINPUT98), .Z(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT99), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT26), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n481), .A2(new_n482), .ZN(new_n729));
  NOR2_X1   g304(.A1(new_n729), .A2(G2105), .ZN(new_n730));
  AOI22_X1  g305(.A1(new_n730), .A2(G141), .B1(G105), .B2(new_n460), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n725), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n723), .B1(new_n733), .B2(new_n708), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT27), .B(G1996), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT88), .B(G16), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G20), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT23), .Z(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G299), .B2(G16), .ZN(new_n740));
  INV_X1    g315(.A(G1956), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n708), .A2(G26), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT28), .Z(new_n744));
  NAND2_X1  g319(.A1(new_n472), .A2(G128), .ZN(new_n745));
  OR2_X1    g320(.A1(G104), .A2(G2105), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n746), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n747));
  INV_X1    g322(.A(G140), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n745), .B(new_n747), .C1(new_n748), .C2(new_n463), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT95), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n744), .B1(new_n751), .B2(G29), .ZN(new_n752));
  INV_X1    g327(.A(G2067), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR4_X1   g329(.A1(new_n722), .A2(new_n736), .A3(new_n742), .A4(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n708), .A2(G33), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n758));
  NAND3_X1  g333(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n730), .A2(G139), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n760), .B(new_n761), .C1(new_n459), .C2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT97), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n757), .B1(new_n764), .B2(G29), .ZN(new_n765));
  INV_X1    g340(.A(G2072), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n720), .A2(new_n721), .ZN(new_n768));
  INV_X1    g343(.A(new_n737), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n769), .A2(G19), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n558), .B2(new_n769), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT94), .B(G1341), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n771), .B(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n708), .A2(G35), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G162), .B2(new_n708), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT29), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n776), .A2(G2090), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n767), .A2(new_n768), .A3(new_n773), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT93), .ZN(new_n779));
  OR3_X1    g354(.A1(new_n779), .A2(G4), .A3(G16), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(G4), .B2(G16), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n605), .A2(new_n608), .ZN(new_n782));
  INV_X1    g357(.A(new_n604), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n780), .B(new_n781), .C1(new_n784), .C2(new_n718), .ZN(new_n785));
  INV_X1    g360(.A(G1348), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n765), .A2(new_n766), .ZN(new_n788));
  NAND2_X1  g363(.A1(G164), .A2(G29), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G27), .B2(G29), .ZN(new_n790));
  INV_X1    g365(.A(G2078), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n776), .A2(G2090), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n790), .A2(new_n791), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n788), .A2(new_n792), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n778), .A2(new_n787), .A3(new_n795), .ZN(new_n796));
  AND3_X1   g371(.A1(new_n706), .A2(new_n755), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT90), .B(KEYINPUT34), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n737), .A2(G22), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G166), .B2(new_n737), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(G1971), .Z(new_n802));
  NAND2_X1  g377(.A1(new_n718), .A2(G23), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n579), .B2(new_n718), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT91), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT33), .B(G1976), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n805), .A2(new_n807), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n802), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n581), .A2(new_n585), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G16), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G6), .B2(G16), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(KEYINPUT32), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n813), .A2(KEYINPUT32), .ZN(new_n816));
  OAI21_X1  g391(.A(G1981), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n816), .ZN(new_n818));
  INV_X1    g393(.A(G1981), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n818), .A2(new_n819), .A3(new_n814), .ZN(new_n820));
  AND2_X1   g395(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n799), .B1(new_n810), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n808), .A2(new_n809), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n817), .A2(new_n820), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n823), .A2(new_n798), .A3(new_n824), .A4(new_n802), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT92), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(KEYINPUT36), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n708), .A2(G25), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n730), .A2(G131), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n472), .A2(G119), .ZN(new_n831));
  OR2_X1    g406(.A1(G95), .A2(G2105), .ZN(new_n832));
  OAI211_X1 g407(.A(new_n832), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n829), .B1(new_n835), .B2(new_n708), .ZN(new_n836));
  XOR2_X1   g411(.A(KEYINPUT35), .B(G1991), .Z(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n836), .B(new_n838), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n737), .A2(G24), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT89), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G290), .B2(new_n769), .ZN(new_n842));
  INV_X1    g417(.A(G1986), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  AOI211_X1 g419(.A(new_n839), .B(new_n844), .C1(new_n826), .C2(KEYINPUT36), .ZN(new_n845));
  NAND4_X1  g420(.A1(new_n822), .A2(new_n825), .A3(new_n828), .A4(new_n845), .ZN(new_n846));
  AND2_X1   g421(.A1(new_n797), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n822), .A2(new_n825), .A3(new_n845), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(new_n827), .ZN(new_n849));
  AND2_X1   g424(.A1(new_n847), .A2(new_n849), .ZN(G311));
  INV_X1    g425(.A(KEYINPUT101), .ZN(new_n851));
  AOI21_X1  g426(.A(new_n851), .B1(new_n847), .B2(new_n849), .ZN(new_n852));
  AND4_X1   g427(.A1(new_n851), .A2(new_n849), .A3(new_n846), .A4(new_n797), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(G150));
  NAND2_X1  g429(.A1(new_n609), .A2(G559), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT38), .Z(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  INV_X1    g432(.A(G67), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n857), .B1(new_n501), .B2(new_n858), .ZN(new_n859));
  AOI22_X1  g434(.A1(new_n859), .A2(G651), .B1(new_n518), .B2(G55), .ZN(new_n860));
  INV_X1    g435(.A(G93), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n861), .B2(new_n526), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n557), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n541), .A2(G93), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n552), .A2(new_n556), .B1(new_n864), .B2(new_n860), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n856), .B(new_n867), .ZN(new_n868));
  AND2_X1   g443(.A1(new_n868), .A2(KEYINPUT39), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n868), .A2(KEYINPUT39), .ZN(new_n870));
  NOR3_X1   g445(.A1(new_n869), .A2(new_n870), .A3(G860), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n862), .A2(G860), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT37), .ZN(new_n873));
  OR2_X1    g448(.A1(new_n871), .A2(new_n873), .ZN(G145));
  XOR2_X1   g449(.A(new_n622), .B(KEYINPUT103), .Z(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n730), .A2(G142), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n877), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT104), .ZN(new_n880));
  OAI21_X1  g455(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n881));
  INV_X1    g456(.A(G118), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n881), .B1(new_n882), .B2(G2105), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(G130), .B2(new_n472), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n879), .A2(new_n880), .A3(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n880), .B1(new_n879), .B2(new_n884), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n886), .A2(new_n835), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n879), .A2(new_n884), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT104), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n834), .B1(new_n890), .B2(new_n885), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n876), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n835), .B1(new_n886), .B2(new_n887), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n834), .A3(new_n885), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n875), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n892), .A2(KEYINPUT105), .A3(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n749), .B(KEYINPUT95), .ZN(new_n897));
  INV_X1    g472(.A(new_n486), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n485), .B1(new_n462), .B2(new_n480), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n472), .A2(G126), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n489), .A2(new_n491), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n897), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n751), .A2(new_n487), .A3(new_n492), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n733), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n904), .A2(new_n905), .A3(new_n733), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n763), .A3(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n764), .ZN(new_n910));
  INV_X1    g485(.A(new_n908), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n910), .B1(new_n911), .B2(new_n906), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n896), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n892), .A2(new_n895), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT105), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n909), .B(new_n912), .C1(new_n915), .C2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(G160), .B(new_n631), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(G162), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n913), .A2(new_n915), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n909), .A2(new_n912), .A3(new_n895), .A4(new_n892), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n919), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g502(.A1(new_n866), .A2(new_n617), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n609), .B(new_n615), .C1(new_n863), .C2(new_n865), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n784), .A2(G299), .ZN(new_n930));
  INV_X1    g505(.A(G299), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n609), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n928), .A2(new_n929), .A3(new_n930), .A4(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT106), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT42), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n928), .A2(new_n929), .ZN(new_n936));
  INV_X1    g511(.A(new_n932), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n609), .A2(new_n931), .ZN(new_n938));
  OAI21_X1  g513(.A(KEYINPUT41), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n930), .A2(new_n940), .A3(new_n932), .ZN(new_n941));
  AOI21_X1  g516(.A(KEYINPUT107), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT107), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n930), .A2(new_n932), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n943), .B1(new_n944), .B2(KEYINPUT41), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n936), .B1(new_n942), .B2(new_n945), .ZN(new_n946));
  AND3_X1   g521(.A1(new_n934), .A2(new_n935), .A3(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n935), .B1(new_n934), .B2(new_n946), .ZN(new_n948));
  XNOR2_X1  g523(.A(G290), .B(G305), .ZN(new_n949));
  XNOR2_X1  g524(.A(G303), .B(G288), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n949), .B(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n951), .ZN(new_n952));
  NOR3_X1   g527(.A1(new_n947), .A2(new_n948), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n934), .A2(new_n946), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT42), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n934), .A2(new_n935), .A3(new_n946), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n951), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(G868), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n862), .A2(new_n595), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(G295));
  INV_X1    g535(.A(KEYINPUT108), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n958), .A2(new_n961), .A3(new_n959), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n952), .B1(new_n947), .B2(new_n948), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n955), .A2(new_n956), .A3(new_n951), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n595), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n959), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT108), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n962), .A2(new_n967), .ZN(G331));
  NAND2_X1  g543(.A1(G171), .A2(KEYINPUT109), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n970));
  NAND2_X1  g545(.A1(G301), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n971), .A3(G286), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n535), .B(new_n536), .ZN(new_n973));
  NAND4_X1  g548(.A1(new_n973), .A2(KEYINPUT109), .A3(new_n531), .A4(G171), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n972), .A2(new_n974), .A3(new_n866), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n972), .A2(new_n974), .A3(KEYINPUT110), .A4(new_n866), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n972), .A2(new_n974), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n944), .B1(new_n980), .B2(new_n867), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n867), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n975), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n939), .A2(new_n941), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n979), .A2(new_n981), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n925), .B1(new_n985), .B2(new_n951), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n981), .A2(new_n975), .ZN(new_n987));
  AOI22_X1  g562(.A1(new_n977), .A2(new_n978), .B1(new_n867), .B2(new_n980), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n942), .A2(new_n945), .ZN(new_n989));
  OAI211_X1 g564(.A(new_n951), .B(new_n987), .C1(new_n988), .C2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT43), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n986), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n987), .B1(new_n988), .B2(new_n989), .ZN(new_n994));
  AOI21_X1  g569(.A(G37), .B1(new_n994), .B2(new_n952), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT43), .B1(new_n995), .B2(new_n990), .ZN(new_n996));
  OAI21_X1  g571(.A(KEYINPUT44), .B1(new_n993), .B2(new_n996), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n986), .A2(new_n991), .A3(KEYINPUT43), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n992), .B1(new_n995), .B2(new_n990), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n997), .B1(new_n1000), .B2(KEYINPUT44), .ZN(G397));
  XNOR2_X1  g576(.A(new_n897), .B(G2067), .ZN(new_n1002));
  INV_X1    g577(.A(G1384), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(new_n900), .B2(new_n903), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT111), .B(KEYINPUT45), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(G125), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n467), .B1(new_n729), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(G2105), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n730), .A2(G137), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(G40), .A4(new_n461), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1006), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1002), .A2(new_n1013), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT113), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n733), .A2(G1996), .ZN(new_n1016));
  INV_X1    g591(.A(G1996), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n732), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1016), .A2(new_n1012), .A3(new_n1018), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(new_n834), .A2(new_n838), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n835), .A2(new_n837), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1012), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1024));
  OR3_X1    g599(.A1(new_n1013), .A2(G290), .A3(G1986), .ZN(new_n1025));
  NAND3_X1  g600(.A1(G290), .A2(G1986), .A3(new_n1012), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1027), .B(KEYINPUT112), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(G40), .ZN(new_n1030));
  NOR3_X1   g605(.A1(new_n465), .A2(new_n468), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT50), .ZN(new_n1032));
  AOI21_X1  g607(.A(G1384), .B1(new_n487), .B2(new_n492), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT66), .B1(new_n900), .B2(new_n903), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n487), .A2(new_n488), .A3(new_n492), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1384), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1034), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g613(.A(KEYINPUT119), .B1(new_n1038), .B2(G1956), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT114), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1005), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1040), .B1(new_n1037), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1003), .B1(new_n493), .B2(new_n494), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(KEYINPUT114), .A3(new_n1005), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1011), .B1(KEYINPUT45), .B2(new_n1033), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT56), .B(G2072), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1043), .A2(KEYINPUT50), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1048), .B(new_n741), .C1(new_n1049), .C2(new_n1034), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1039), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT122), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT57), .ZN(new_n1054));
  AND3_X1   g629(.A1(G299), .A2(KEYINPUT120), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(KEYINPUT120), .B1(G299), .B2(new_n1054), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND4_X1  g632(.A1(new_n568), .A2(new_n569), .A3(KEYINPUT57), .A4(new_n573), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT121), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1057), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1039), .A2(new_n1047), .A3(new_n1050), .A4(KEYINPUT122), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1053), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1060), .A2(new_n1039), .A3(new_n1047), .A4(new_n1050), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1064), .A2(KEYINPUT61), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT61), .ZN(new_n1067));
  AND2_X1   g642(.A1(new_n1051), .A2(new_n1061), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1064), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1011), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1071), .B1(new_n1037), .B2(new_n1032), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n786), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1031), .A2(new_n753), .A3(new_n1033), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT60), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1032), .B(new_n1003), .C1(new_n900), .C2(new_n903), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1076), .A2(new_n1031), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1077), .B1(new_n1043), .B2(KEYINPUT50), .ZN(new_n1078));
  OAI211_X1 g653(.A(KEYINPUT60), .B(new_n1074), .C1(new_n1078), .C2(G1348), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n609), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1073), .A2(KEYINPUT60), .A3(new_n784), .A4(new_n1074), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1075), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1042), .A2(new_n1017), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1084));
  XOR2_X1   g659(.A(KEYINPUT58), .B(G1341), .Z(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(new_n558), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT59), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1087), .A2(new_n1090), .A3(new_n558), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1082), .B1(new_n1089), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1066), .A2(new_n1070), .A3(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n784), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1064), .A2(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1063), .A2(new_n1095), .ZN(new_n1096));
  AND3_X1   g671(.A1(new_n1093), .A2(KEYINPUT123), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT123), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1042), .A2(new_n791), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT45), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1011), .B1(new_n1004), .B2(new_n1102), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1100), .A2(G2078), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1103), .B(new_n1104), .C1(new_n1043), .C2(new_n1005), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1072), .A2(new_n721), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1101), .A2(G301), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1011), .A2(KEYINPUT125), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1033), .A2(KEYINPUT45), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1011), .A2(KEYINPUT125), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1006), .A2(new_n1104), .ZN(new_n1112));
  NOR2_X1   g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI221_X4 g688(.A(new_n1113), .B1(new_n721), .B2(new_n1072), .C1(new_n1099), .C2(new_n1100), .ZN(new_n1114));
  OAI211_X1 g689(.A(KEYINPUT54), .B(new_n1107), .C1(new_n1114), .C2(G301), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1103), .B1(new_n1043), .B2(new_n1005), .ZN(new_n1117));
  INV_X1    g692(.A(G1966), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1119), .B1(G2084), .B2(new_n1072), .ZN(new_n1120));
  OAI211_X1 g695(.A(new_n1116), .B(G8), .C1(new_n1120), .C2(G286), .ZN(new_n1121));
  NAND2_X1  g696(.A1(G286), .A2(G8), .ZN(new_n1122));
  INV_X1    g697(.A(G2084), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1123), .A2(new_n1078), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1124));
  INV_X1    g699(.A(G8), .ZN(new_n1125));
  OAI211_X1 g700(.A(KEYINPUT51), .B(new_n1122), .C1(new_n1124), .C2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1122), .ZN(new_n1127));
  AOI21_X1  g702(.A(KEYINPUT124), .B1(new_n1120), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1124), .A2(new_n1129), .A3(new_n1122), .ZN(new_n1130));
  OAI211_X1 g705(.A(new_n1121), .B(new_n1126), .C1(new_n1128), .C2(new_n1130), .ZN(new_n1131));
  AND2_X1   g706(.A1(new_n1115), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n521), .A2(new_n527), .A3(G8), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n1133), .B(KEYINPUT55), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1042), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1135));
  XNOR2_X1  g710(.A(KEYINPUT115), .B(G1971), .ZN(new_n1136));
  INV_X1    g711(.A(G2090), .ZN(new_n1137));
  AOI22_X1  g712(.A1(new_n1135), .A2(new_n1136), .B1(new_n1137), .B2(new_n1038), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1134), .B1(new_n1138), .B2(new_n1125), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1084), .A2(G8), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n811), .A2(new_n819), .ZN(new_n1141));
  NAND2_X1  g716(.A1(G305), .A2(G1981), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT49), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1140), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1144), .B2(new_n1143), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1140), .B1(G1976), .B2(new_n579), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT52), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1147), .B(new_n1148), .C1(G1976), .C2(new_n579), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1146), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1152));
  AOI21_X1  g727(.A(KEYINPUT114), .B1(new_n1043), .B2(new_n1005), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1136), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1137), .B(new_n1071), .C1(new_n1037), .C2(new_n1032), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1134), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1156), .A2(G8), .A3(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT116), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1125), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1161), .A2(KEYINPUT116), .A3(new_n1157), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1151), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT54), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1101), .A2(new_n1106), .ZN(new_n1165));
  NOR3_X1   g740(.A1(new_n1165), .A2(G171), .A3(new_n1113), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1099), .A2(new_n1100), .B1(new_n721), .B2(new_n1072), .ZN(new_n1167));
  AOI21_X1  g742(.A(G301), .B1(new_n1167), .B2(new_n1105), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1164), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1132), .A2(new_n1139), .A3(new_n1163), .A4(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1097), .A2(new_n1098), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT118), .ZN(new_n1172));
  AOI21_X1  g747(.A(KEYINPUT116), .B1(new_n1161), .B2(new_n1157), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1155), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1174), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1175));
  NOR4_X1   g750(.A1(new_n1175), .A2(new_n1159), .A3(new_n1125), .A4(new_n1134), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1173), .A2(new_n1176), .A3(new_n1151), .ZN(new_n1177));
  INV_X1    g752(.A(G1976), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1146), .A2(new_n1178), .A3(new_n579), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1141), .B(KEYINPUT117), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1140), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1172), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1181), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1146), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1184));
  NAND3_X1  g759(.A1(new_n1160), .A2(new_n1162), .A3(new_n1184), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1183), .A2(new_n1185), .A3(KEYINPUT118), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1182), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n1188));
  OAI211_X1 g763(.A(new_n1139), .B(new_n1184), .C1(new_n1173), .C2(new_n1176), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1120), .A2(G8), .A3(G168), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NOR2_X1   g766(.A1(new_n1161), .A2(new_n1157), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1192), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1163), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1191), .A2(new_n1194), .ZN(new_n1195));
  OR2_X1    g770(.A1(new_n1131), .A2(KEYINPUT62), .ZN(new_n1196));
  INV_X1    g771(.A(new_n1168), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1197), .B1(new_n1131), .B2(KEYINPUT62), .ZN(new_n1198));
  NAND4_X1  g773(.A1(new_n1196), .A2(new_n1198), .A3(new_n1139), .A4(new_n1163), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1187), .A2(new_n1195), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1029), .B1(new_n1171), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1012), .A2(new_n1017), .ZN(new_n1202));
  INV_X1    g777(.A(KEYINPUT46), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  XOR2_X1   g779(.A(new_n1204), .B(KEYINPUT126), .Z(new_n1205));
  AOI21_X1  g780(.A(new_n1013), .B1(new_n1002), .B2(new_n733), .ZN(new_n1206));
  AOI21_X1  g781(.A(new_n1206), .B1(new_n1203), .B2(new_n1202), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT47), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1025), .B(KEYINPUT48), .Z(new_n1210));
  OAI21_X1  g785(.A(new_n1209), .B1(new_n1024), .B2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1212));
  NAND2_X1  g787(.A1(new_n897), .A2(new_n753), .ZN(new_n1213));
  AOI21_X1  g788(.A(new_n1013), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1201), .A2(new_n1215), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g791(.A1(new_n994), .A2(new_n952), .ZN(new_n1218));
  NAND3_X1  g792(.A1(new_n1218), .A2(new_n925), .A3(new_n990), .ZN(new_n1219));
  NAND2_X1  g793(.A1(new_n1219), .A2(KEYINPUT43), .ZN(new_n1220));
  OR2_X1    g794(.A1(new_n985), .A2(new_n951), .ZN(new_n1221));
  NAND4_X1  g795(.A1(new_n1221), .A2(new_n992), .A3(new_n925), .A4(new_n990), .ZN(new_n1222));
  NAND2_X1  g796(.A1(new_n1220), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g797(.A1(new_n669), .A2(G319), .A3(new_n650), .ZN(new_n1224));
  NOR2_X1   g798(.A1(new_n1224), .A2(G229), .ZN(new_n1225));
  NAND2_X1  g799(.A1(new_n926), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g800(.A(new_n1226), .ZN(new_n1227));
  AOI21_X1  g801(.A(KEYINPUT127), .B1(new_n1223), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n1229));
  AOI211_X1 g803(.A(new_n1229), .B(new_n1226), .C1(new_n1220), .C2(new_n1222), .ZN(new_n1230));
  NOR2_X1   g804(.A1(new_n1228), .A2(new_n1230), .ZN(G308));
  OAI21_X1  g805(.A(new_n1229), .B1(new_n1000), .B2(new_n1226), .ZN(new_n1232));
  NAND3_X1  g806(.A1(new_n1223), .A2(KEYINPUT127), .A3(new_n1227), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n1232), .A2(new_n1233), .ZN(G225));
endmodule


