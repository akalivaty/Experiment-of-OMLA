//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n210));
  NAND2_X1  g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n208), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  OR2_X1    g0015(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n208), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT0), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n204), .A2(new_n205), .ZN(new_n220));
  INV_X1    g0020(.A(G50), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G1), .A2(G13), .ZN(new_n223));
  INV_X1    g0023(.A(G20), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n222), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n216), .A2(new_n219), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n215), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G50), .B(G68), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT65), .ZN(new_n239));
  XOR2_X1   g0039(.A(G58), .B(G77), .Z(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(KEYINPUT66), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n241), .B(new_n245), .Z(G351));
  OR2_X1    g0046(.A1(KEYINPUT3), .A2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(KEYINPUT3), .A2(G33), .ZN(new_n248));
  AOI21_X1  g0048(.A(G1698), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(G222), .ZN(new_n250));
  INV_X1    g0050(.A(G77), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT3), .B(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G223), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(G1698), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n250), .B1(new_n251), .B2(new_n252), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  AND2_X1   g0055(.A1(G33), .A2(G41), .ZN(new_n256));
  NOR3_X1   g0056(.A1(new_n256), .A2(KEYINPUT67), .A3(new_n223), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT67), .ZN(new_n258));
  AND2_X1   g0058(.A1(G1), .A2(G13), .ZN(new_n259));
  NAND2_X1  g0059(.A1(G33), .A2(G41), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n257), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  AOI21_X1  g0065(.A(G1), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n260), .A2(G1), .A3(G13), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(new_n267), .A3(G274), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G1), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n270), .B1(G41), .B2(G45), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n269), .B1(G226), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n263), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G190), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G200), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n278), .B1(new_n263), .B2(new_n274), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n270), .A2(G13), .A3(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n221), .ZN(new_n282));
  INV_X1    g0082(.A(new_n281), .ZN(new_n283));
  NAND3_X1  g0083(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n223), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT69), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT69), .B1(new_n283), .B2(new_n285), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n288), .A2(new_n289), .B1(new_n270), .B2(G20), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n282), .B1(new_n290), .B2(new_n221), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT70), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XOR2_X1   g0093(.A(KEYINPUT8), .B(G58), .Z(new_n294));
  NOR2_X1   g0094(.A1(new_n294), .A2(KEYINPUT68), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT68), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n296), .A2(new_n202), .A3(KEYINPUT8), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n224), .A2(G33), .ZN(new_n300));
  INV_X1    g0100(.A(G150), .ZN(new_n301));
  INV_X1    g0101(.A(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n224), .A2(new_n302), .ZN(new_n303));
  OAI22_X1  g0103(.A1(new_n299), .A2(new_n300), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n224), .B1(new_n220), .B2(new_n221), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n285), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n293), .A2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n307), .A2(KEYINPUT9), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n309), .B1(new_n293), .B2(new_n306), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n280), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT10), .B1(new_n279), .B2(KEYINPUT72), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g0114(.A(new_n312), .B(new_n280), .C1(new_n308), .C2(new_n310), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n275), .A2(G179), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n317), .B1(new_n318), .B2(new_n275), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n307), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT71), .ZN(new_n322));
  NOR2_X1   g0122(.A1(G20), .A2(G33), .ZN(new_n323));
  AOI22_X1  g0123(.A1(new_n294), .A2(new_n323), .B1(G20), .B2(G77), .ZN(new_n324));
  XNOR2_X1  g0124(.A(KEYINPUT15), .B(G87), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n324), .B1(new_n300), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n285), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n251), .B1(new_n270), .B2(G20), .ZN(new_n328));
  AOI22_X1  g0128(.A1(new_n286), .A2(new_n328), .B1(new_n251), .B2(new_n283), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n249), .A2(G232), .ZN(new_n331));
  INV_X1    g0131(.A(G107), .ZN(new_n332));
  INV_X1    g0132(.A(G238), .ZN(new_n333));
  OAI221_X1 g0133(.A(new_n331), .B1(new_n332), .B2(new_n252), .C1(new_n333), .C2(new_n254), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n262), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n269), .B1(G244), .B2(new_n273), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n322), .B(new_n330), .C1(new_n337), .C2(G169), .ZN(new_n338));
  AOI21_X1  g0138(.A(G169), .B1(new_n335), .B2(new_n336), .ZN(new_n339));
  INV_X1    g0139(.A(new_n330), .ZN(new_n340));
  OAI21_X1  g0140(.A(KEYINPUT71), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(G179), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n337), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n338), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n330), .B1(new_n337), .B2(G190), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n345), .B1(new_n278), .B2(new_n337), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT13), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT73), .ZN(new_n349));
  INV_X1    g0149(.A(G97), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n302), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g0151(.A1(G226), .A2(G1698), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(new_n230), .B2(G1698), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n351), .B1(new_n353), .B2(new_n252), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n267), .A2(KEYINPUT67), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n259), .A2(new_n258), .A3(new_n260), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n349), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n230), .A2(G1698), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n359), .B1(G226), .B2(G1698), .ZN(new_n360));
  AND2_X1   g0160(.A1(KEYINPUT3), .A2(G33), .ZN(new_n361));
  NOR2_X1   g0161(.A1(KEYINPUT3), .A2(G33), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n360), .A2(new_n363), .B1(new_n302), .B2(new_n350), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(new_n262), .A3(KEYINPUT73), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n358), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n268), .B1(new_n333), .B2(new_n272), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n348), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  AOI211_X1 g0169(.A(KEYINPUT13), .B(new_n367), .C1(new_n358), .C2(new_n365), .ZN(new_n370));
  OAI21_X1  g0170(.A(G169), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(KEYINPUT14), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n366), .A2(new_n368), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT74), .B1(new_n373), .B2(KEYINPUT13), .ZN(new_n374));
  INV_X1    g0174(.A(new_n369), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT74), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n366), .A2(new_n376), .A3(new_n348), .A4(new_n368), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n374), .A2(new_n375), .A3(G179), .A4(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT14), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n379), .B(G169), .C1(new_n369), .C2(new_n370), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n372), .A2(new_n378), .A3(new_n380), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n284), .A2(new_n223), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n323), .A2(G50), .ZN(new_n383));
  XOR2_X1   g0183(.A(new_n383), .B(KEYINPUT75), .Z(new_n384));
  OAI22_X1  g0184(.A1(new_n300), .A2(new_n251), .B1(new_n224), .B2(G68), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n382), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n387), .A2(KEYINPUT11), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(KEYINPUT11), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT12), .B1(new_n281), .B2(G68), .ZN(new_n390));
  OR3_X1    g0190(.A1(new_n281), .A2(KEYINPUT12), .A3(G68), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n203), .B1(new_n270), .B2(G20), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n390), .A2(new_n391), .B1(new_n286), .B2(new_n392), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n381), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n374), .A2(new_n375), .A3(G190), .A4(new_n377), .ZN(new_n396));
  INV_X1    g0196(.A(new_n394), .ZN(new_n397));
  OAI21_X1  g0197(.A(G200), .B1(new_n369), .B2(new_n370), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n347), .A2(new_n395), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT16), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT7), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n252), .B2(G20), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n363), .A2(KEYINPUT7), .A3(new_n224), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n401), .B1(new_n405), .B2(G68), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G58), .A2(G68), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n204), .A2(new_n205), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G20), .ZN(new_n409));
  INV_X1    g0209(.A(G159), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n303), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT76), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT76), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n409), .A2(new_n415), .A3(new_n412), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n406), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n203), .B1(new_n403), .B2(new_n404), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n401), .B1(new_n418), .B2(new_n413), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n285), .A3(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n298), .A2(new_n283), .ZN(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n290), .B2(new_n299), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G1698), .ZN(new_n425));
  OAI211_X1 g0225(.A(G223), .B(new_n425), .C1(new_n361), .C2(new_n362), .ZN(new_n426));
  OAI211_X1 g0226(.A(G226), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G87), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n357), .B1(new_n429), .B2(KEYINPUT77), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT77), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n426), .A2(new_n427), .A3(new_n431), .A4(new_n428), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n268), .B1(new_n230), .B2(new_n272), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT78), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT78), .ZN(new_n436));
  OAI211_X1 g0236(.A(new_n268), .B(new_n436), .C1(new_n230), .C2(new_n272), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n433), .A2(new_n438), .A3(G179), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n430), .A2(new_n432), .B1(new_n435), .B2(new_n437), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(new_n318), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n424), .A2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(KEYINPUT18), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n433), .A2(new_n438), .A3(new_n276), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(G200), .B1(new_n433), .B2(new_n438), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n420), .B(new_n423), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT17), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT18), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n424), .A2(new_n450), .A3(new_n441), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n444), .B1(G200), .B2(new_n440), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n452), .A2(KEYINPUT17), .A3(new_n420), .A4(new_n423), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n443), .A2(new_n449), .A3(new_n451), .A4(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n400), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n321), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(G264), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n457));
  OAI211_X1 g0257(.A(G257), .B(new_n425), .C1(new_n361), .C2(new_n362), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n247), .A2(G303), .A3(new_n248), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT87), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n457), .A2(new_n458), .A3(KEYINPUT87), .A4(new_n459), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n262), .A3(new_n463), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n270), .B(G45), .C1(new_n264), .C2(KEYINPUT5), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT79), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n265), .A2(G1), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT79), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT5), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(G41), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n467), .A2(new_n468), .A3(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(G274), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(new_n259), .B2(new_n260), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n469), .A2(G41), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n466), .A2(new_n471), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  OAI211_X1 g0276(.A(G270), .B(new_n267), .C1(new_n465), .C2(new_n474), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT86), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT86), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n480), .A3(new_n477), .ZN(new_n481));
  AND3_X1   g0281(.A1(new_n464), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(G33), .A2(G283), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n483), .B(new_n224), .C1(G33), .C2(new_n350), .ZN(new_n484));
  INV_X1    g0284(.A(G116), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n485), .A2(G20), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n285), .A3(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT20), .ZN(new_n488));
  XNOR2_X1  g0288(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n281), .A2(G116), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n270), .A2(G33), .ZN(new_n491));
  AND3_X1   g0291(.A1(new_n382), .A2(new_n281), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n490), .B1(new_n492), .B2(G116), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n482), .A2(new_n494), .A3(G179), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n464), .A2(new_n479), .A3(new_n481), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT21), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n318), .B1(new_n489), .B2(new_n493), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n496), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n497), .B1(new_n496), .B2(new_n498), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n495), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n482), .A2(G190), .ZN(new_n502));
  INV_X1    g0302(.A(new_n494), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n496), .A2(G200), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT88), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT88), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n502), .A2(new_n507), .A3(new_n503), .A4(new_n504), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n501), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n332), .A2(G20), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT90), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT23), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n224), .A2(G33), .A3(G116), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n510), .B2(KEYINPUT23), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n511), .B1(new_n510), .B2(KEYINPUT23), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n224), .B(G87), .C1(new_n361), .C2(new_n362), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT22), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT22), .ZN(new_n520));
  NAND4_X1  g0320(.A1(new_n252), .A2(new_n520), .A3(new_n224), .A4(G87), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT91), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n517), .A2(new_n522), .A3(KEYINPUT91), .ZN(new_n526));
  XNOR2_X1  g0326(.A(KEYINPUT89), .B(KEYINPUT24), .ZN(new_n527));
  INV_X1    g0327(.A(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n525), .A2(new_n526), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g0329(.A(KEYINPUT91), .B1(new_n517), .B2(new_n522), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n382), .B1(new_n530), .B2(new_n527), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT25), .B1(new_n283), .B2(new_n332), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n283), .A2(KEYINPUT25), .A3(new_n332), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n534), .A2(new_n535), .B1(new_n492), .B2(G107), .ZN(new_n536));
  OAI211_X1 g0336(.A(G257), .B(G1698), .C1(new_n361), .C2(new_n362), .ZN(new_n537));
  OAI211_X1 g0337(.A(G250), .B(new_n425), .C1(new_n361), .C2(new_n362), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G33), .A2(G294), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n262), .ZN(new_n541));
  OAI211_X1 g0341(.A(G264), .B(new_n267), .C1(new_n465), .C2(new_n474), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n541), .A2(new_n476), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(new_n278), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(G190), .B2(new_n543), .ZN(new_n545));
  AND3_X1   g0345(.A1(new_n532), .A2(new_n536), .A3(new_n545), .ZN(new_n546));
  AND3_X1   g0346(.A1(new_n541), .A2(G179), .A3(new_n542), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(new_n476), .B1(new_n543), .B2(G169), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n548), .B1(new_n532), .B2(new_n536), .ZN(new_n549));
  OAI21_X1  g0349(.A(KEYINPUT92), .B1(new_n546), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n536), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n529), .B2(new_n531), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n545), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT92), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n553), .B(new_n554), .C1(new_n552), .C2(new_n548), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n249), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n252), .A2(G244), .A3(G1698), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n357), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n267), .A2(G274), .A3(new_n467), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT82), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n473), .A2(KEYINPUT82), .A3(new_n467), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n256), .A2(new_n223), .ZN(new_n566));
  OAI21_X1  g0366(.A(G250), .B1(new_n265), .B2(G1), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(KEYINPUT83), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT83), .ZN(new_n571));
  AOI211_X1 g0371(.A(new_n571), .B(new_n568), .C1(new_n563), .C2(new_n564), .ZN(new_n572));
  OAI211_X1 g0372(.A(G179), .B(new_n560), .C1(new_n570), .C2(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT82), .B1(new_n473), .B2(new_n467), .ZN(new_n574));
  AND4_X1   g0374(.A1(KEYINPUT82), .A2(new_n267), .A3(G274), .A4(new_n467), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n569), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n571), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n565), .A2(KEYINPUT83), .A3(new_n569), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n559), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n573), .B1(new_n579), .B2(new_n318), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT84), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n573), .B(KEYINPUT84), .C1(new_n579), .C2(new_n318), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n252), .A2(new_n224), .A3(G68), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n300), .B2(new_n350), .ZN(new_n586));
  XNOR2_X1  g0386(.A(KEYINPUT85), .B(G87), .ZN(new_n587));
  NOR2_X1   g0387(.A1(G97), .A2(G107), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(G20), .B1(new_n351), .B2(KEYINPUT19), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n584), .B(new_n586), .C1(new_n590), .C2(new_n591), .ZN(new_n592));
  AOI22_X1  g0392(.A1(new_n592), .A2(new_n285), .B1(new_n283), .B2(new_n325), .ZN(new_n593));
  INV_X1    g0393(.A(new_n492), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n325), .B2(new_n594), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n582), .A2(new_n583), .A3(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT80), .ZN(new_n597));
  OAI211_X1 g0397(.A(G257), .B(new_n267), .C1(new_n465), .C2(new_n474), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n476), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n597), .B1(new_n476), .B2(new_n598), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g0401(.A(G244), .B(new_n425), .C1(new_n361), .C2(new_n362), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT4), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n252), .A2(KEYINPUT4), .A3(G244), .A4(new_n425), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n252), .A2(G250), .A3(G1698), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n483), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n607), .A2(new_n262), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n601), .A2(KEYINPUT81), .A3(new_n342), .A4(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n281), .A2(G97), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n492), .B2(G97), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n332), .A2(KEYINPUT6), .A3(G97), .ZN(new_n613));
  XOR2_X1   g0413(.A(G97), .B(G107), .Z(new_n614));
  OAI21_X1  g0414(.A(new_n613), .B1(new_n614), .B2(KEYINPUT6), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n615), .A2(G20), .B1(G77), .B2(new_n323), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n405), .A2(G107), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n612), .B1(new_n618), .B2(new_n285), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT81), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n476), .A2(new_n598), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(KEYINPUT80), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n476), .A2(new_n597), .A3(new_n598), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n623), .A2(new_n608), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n621), .B1(new_n625), .B2(new_n318), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(G179), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n609), .B(new_n620), .C1(new_n626), .C2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n577), .A2(new_n578), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(G190), .A3(new_n560), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n492), .A2(G87), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n593), .A2(new_n631), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n630), .B(new_n632), .C1(new_n278), .C2(new_n579), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n625), .A2(G200), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n634), .B(new_n619), .C1(new_n276), .C2(new_n625), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n628), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n596), .A2(new_n636), .ZN(new_n637));
  AND4_X1   g0437(.A1(new_n456), .A2(new_n509), .A3(new_n556), .A4(new_n637), .ZN(G372));
  NAND2_X1  g0438(.A1(new_n449), .A2(new_n453), .ZN(new_n639));
  INV_X1    g0439(.A(new_n344), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n399), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n639), .B1(new_n641), .B2(new_n395), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n443), .A2(new_n451), .ZN(new_n643));
  INV_X1    g0443(.A(new_n643), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n316), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n320), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n456), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n580), .A2(new_n595), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n628), .A2(new_n633), .A3(new_n553), .A4(new_n635), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n501), .A2(new_n549), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT26), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n649), .A2(new_n633), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n653), .B1(new_n654), .B2(new_n628), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n582), .A2(new_n583), .A3(new_n595), .ZN(new_n656));
  INV_X1    g0456(.A(new_n628), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n656), .A2(KEYINPUT26), .A3(new_n657), .A4(new_n633), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n652), .B1(new_n655), .B2(new_n658), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n647), .B1(new_n648), .B2(new_n659), .ZN(G369));
  NAND3_X1  g0460(.A1(new_n270), .A2(new_n224), .A3(G13), .ZN(new_n661));
  OR2_X1    g0461(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(KEYINPUT27), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(G213), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(G343), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n503), .A2(new_n667), .ZN(new_n668));
  MUX2_X1   g0468(.A(new_n509), .B(new_n501), .S(new_n668), .Z(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G330), .ZN(new_n670));
  INV_X1    g0470(.A(new_n552), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n666), .ZN(new_n672));
  AOI22_X1  g0472(.A1(new_n556), .A2(new_n672), .B1(new_n549), .B2(new_n666), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n556), .A2(new_n501), .A3(new_n667), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n549), .A2(new_n667), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n217), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n589), .A2(G116), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(new_n683), .A3(G1), .ZN(new_n684));
  INV_X1    g0484(.A(new_n222), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(new_n682), .ZN(new_n686));
  XNOR2_X1  g0486(.A(new_n686), .B(KEYINPUT28), .ZN(new_n687));
  INV_X1    g0487(.A(new_n649), .ZN(new_n688));
  INV_X1    g0488(.A(new_n650), .ZN(new_n689));
  INV_X1    g0489(.A(new_n651), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n658), .A2(new_n655), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n693), .A2(new_n667), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(KEYINPUT29), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n656), .A2(new_n653), .A3(new_n657), .A4(new_n633), .ZN(new_n696));
  OAI21_X1  g0496(.A(KEYINPUT26), .B1(new_n654), .B2(new_n628), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n667), .B1(new_n698), .B2(new_n652), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n699), .A2(KEYINPUT29), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n695), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G330), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n637), .A2(new_n509), .A3(new_n556), .A4(new_n667), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n623), .A2(new_n608), .A3(new_n624), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n482), .A2(new_n705), .A3(new_n579), .A4(new_n547), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n476), .A2(new_n480), .A3(new_n477), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n480), .B1(new_n476), .B2(new_n477), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n629), .A2(new_n560), .B1(new_n710), .B2(new_n464), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n543), .A2(new_n342), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n712), .B1(new_n608), .B2(new_n601), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n706), .A2(new_n707), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  AND3_X1   g0514(.A1(new_n601), .A2(new_n547), .A3(new_n608), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n715), .A2(KEYINPUT30), .A3(new_n482), .A4(new_n579), .ZN(new_n716));
  AOI211_X1 g0516(.A(new_n704), .B(new_n667), .C1(new_n714), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n706), .A2(new_n707), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n711), .A2(new_n713), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(new_n716), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(KEYINPUT31), .B1(new_n720), .B2(new_n666), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n717), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n702), .B1(new_n703), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n701), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n687), .B1(new_n726), .B2(G1), .ZN(G364));
  INV_X1    g0527(.A(G13), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G20), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n270), .B1(new_n729), .B2(G45), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n681), .A2(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n669), .B2(G330), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G330), .B2(new_n669), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n680), .A2(new_n363), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G355), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G116), .B2(new_n217), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n241), .A2(G45), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n680), .A2(new_n252), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n740), .B1(new_n222), .B2(new_n265), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n737), .B1(new_n738), .B2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n224), .B1(KEYINPUT93), .B2(new_n318), .ZN(new_n743));
  OR2_X1    g0543(.A1(new_n318), .A2(KEYINPUT93), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n223), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(G13), .A2(G33), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G20), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n732), .B1(new_n742), .B2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(G20), .A2(G179), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT94), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n276), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n221), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n224), .A2(G179), .ZN(new_n758));
  NOR2_X1   g0558(.A1(G190), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G159), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n762), .B(KEYINPUT32), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n758), .A2(G190), .A3(G200), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n252), .B1(new_n764), .B2(new_n587), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n276), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n766), .A2(new_n342), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G20), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n758), .A2(new_n276), .A3(G200), .ZN(new_n770));
  OAI22_X1  g0570(.A1(new_n769), .A2(new_n350), .B1(new_n770), .B2(new_n332), .ZN(new_n771));
  NOR4_X1   g0571(.A1(new_n757), .A2(new_n763), .A3(new_n765), .A4(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n753), .A2(new_n766), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n753), .A2(new_n759), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n202), .A2(new_n773), .B1(new_n774), .B2(new_n251), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT95), .Z(new_n776));
  NAND3_X1  g0576(.A1(new_n753), .A2(new_n276), .A3(G200), .ZN(new_n777));
  INV_X1    g0577(.A(KEYINPUT96), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n777), .A2(new_n778), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n772), .B(new_n776), .C1(new_n203), .C2(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G311), .ZN(new_n784));
  INV_X1    g0584(.A(G322), .ZN(new_n785));
  OAI22_X1  g0585(.A1(new_n784), .A2(new_n774), .B1(new_n773), .B2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(G294), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n769), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(G329), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n363), .B1(new_n760), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(G283), .ZN(new_n791));
  INV_X1    g0591(.A(G303), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(new_n770), .B1(new_n764), .B2(new_n792), .ZN(new_n793));
  NOR4_X1   g0593(.A1(new_n786), .A2(new_n788), .A3(new_n790), .A4(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(G326), .ZN(new_n795));
  XOR2_X1   g0595(.A(KEYINPUT33), .B(G317), .Z(new_n796));
  OAI221_X1 g0596(.A(new_n794), .B1(new_n795), .B2(new_n756), .C1(new_n782), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n783), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n751), .B1(new_n798), .B2(new_n745), .ZN(new_n799));
  INV_X1    g0599(.A(new_n748), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n799), .B1(new_n669), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g0601(.A1(new_n734), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  INV_X1    g0603(.A(KEYINPUT98), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n347), .A2(new_n667), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n659), .B2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n805), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n693), .A2(KEYINPUT98), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n694), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n340), .A2(new_n667), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n344), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n812), .B1(new_n347), .B2(new_n811), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n809), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n732), .B1(new_n815), .B2(new_n724), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n816), .B1(new_n724), .B2(new_n815), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n745), .A2(new_n746), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n363), .B1(new_n760), .B2(new_n784), .ZN(new_n820));
  INV_X1    g0620(.A(G87), .ZN(new_n821));
  OAI22_X1  g0621(.A1(new_n821), .A2(new_n770), .B1(new_n764), .B2(new_n332), .ZN(new_n822));
  AOI211_X1 g0622(.A(new_n820), .B(new_n822), .C1(G97), .C2(new_n768), .ZN(new_n823));
  INV_X1    g0623(.A(new_n774), .ZN(new_n824));
  INV_X1    g0624(.A(new_n773), .ZN(new_n825));
  AOI22_X1  g0625(.A1(G116), .A2(new_n824), .B1(new_n825), .B2(G294), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n823), .B(new_n826), .C1(new_n792), .C2(new_n756), .ZN(new_n827));
  INV_X1    g0627(.A(new_n782), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n827), .B1(new_n828), .B2(G283), .ZN(new_n829));
  AOI22_X1  g0629(.A1(G143), .A2(new_n825), .B1(new_n824), .B2(G159), .ZN(new_n830));
  INV_X1    g0630(.A(G137), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n830), .B1(new_n831), .B2(new_n756), .C1(new_n782), .C2(new_n301), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT34), .ZN(new_n833));
  INV_X1    g0633(.A(G132), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n252), .B1(new_n760), .B2(new_n834), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n769), .A2(new_n202), .B1(new_n764), .B2(new_n221), .ZN(new_n836));
  INV_X1    g0636(.A(new_n770), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n835), .B(new_n836), .C1(G68), .C2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n829), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n745), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n732), .B1(G77), .B2(new_n819), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  XOR2_X1   g0641(.A(new_n841), .B(KEYINPUT97), .Z(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n747), .B2(new_n814), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n817), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G384));
  NOR2_X1   g0645(.A1(new_n729), .A2(new_n270), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT103), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT101), .ZN(new_n848));
  INV_X1    g0648(.A(new_n290), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n421), .B1(new_n849), .B2(new_n298), .ZN(new_n850));
  AOI211_X1 g0650(.A(KEYINPUT76), .B(new_n411), .C1(new_n408), .C2(G20), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n415), .B1(new_n409), .B2(new_n412), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n382), .B1(new_n853), .B2(new_n406), .ZN(new_n854));
  INV_X1    g0654(.A(new_n418), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n855), .A2(new_n414), .A3(new_n416), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n401), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n850), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n848), .B1(new_n858), .B2(new_n664), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n417), .A2(new_n285), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT16), .B1(new_n853), .B2(new_n855), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n423), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n664), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n862), .A2(KEYINPUT101), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n454), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n424), .A2(new_n863), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT37), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n442), .A2(new_n868), .A3(new_n869), .A4(new_n447), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n862), .A2(new_n441), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n859), .A2(new_n864), .A3(new_n447), .A4(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n871), .B1(KEYINPUT37), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n847), .B1(new_n867), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n870), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n877), .A2(KEYINPUT103), .A3(KEYINPUT38), .A4(new_n866), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n442), .A2(new_n868), .A3(new_n447), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n880), .A2(KEYINPUT37), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n870), .ZN(new_n882));
  INV_X1    g0682(.A(new_n868), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n882), .A2(KEYINPUT102), .B1(new_n454), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT102), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n881), .A2(new_n885), .A3(new_n870), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT38), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  OAI21_X1  g0687(.A(KEYINPUT105), .B1(new_n879), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n882), .A2(KEYINPUT102), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n454), .A2(new_n883), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(new_n886), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT105), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n893), .A2(new_n894), .A3(new_n875), .A4(new_n878), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n703), .A2(new_n722), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n394), .A2(new_n666), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT100), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n395), .A2(new_n898), .A3(new_n399), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n395), .A2(KEYINPUT100), .A3(new_n399), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n901), .A2(new_n381), .A3(new_n897), .ZN(new_n902));
  AOI22_X1  g0702(.A1(new_n897), .A2(new_n899), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n896), .A2(new_n903), .A3(new_n814), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT40), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n888), .A2(new_n895), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(KEYINPUT106), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT106), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n888), .A2(new_n906), .A3(new_n895), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n908), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n454), .A2(new_n865), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n892), .B1(new_n874), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n877), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n914));
  AND2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n905), .B1(new_n915), .B2(new_n904), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n911), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT107), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n456), .A2(new_n896), .ZN(new_n919));
  INV_X1    g0719(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n702), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n918), .B2(new_n920), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT39), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n879), .B2(new_n887), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT39), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n395), .A2(new_n666), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n644), .A2(new_n664), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n640), .A2(new_n667), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT98), .B1(new_n693), .B2(new_n807), .ZN(new_n931));
  AOI211_X1 g0731(.A(new_n804), .B(new_n805), .C1(new_n691), .C2(new_n692), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n930), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n915), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n933), .A2(new_n934), .A3(new_n903), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n928), .A2(new_n929), .A3(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(KEYINPUT104), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(new_n903), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(new_n809), .B2(new_n930), .ZN(new_n940));
  AOI22_X1  g0740(.A1(new_n940), .A2(new_n934), .B1(new_n644), .B2(new_n664), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(KEYINPUT104), .A3(new_n928), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n938), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n701), .A2(new_n648), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n944), .A2(new_n646), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n943), .B(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n846), .B1(new_n922), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n946), .B2(new_n922), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n615), .A2(KEYINPUT35), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n615), .A2(KEYINPUT35), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n949), .A2(G116), .A3(new_n225), .A4(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT36), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n222), .A2(G77), .A3(new_n407), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(G50), .B2(new_n203), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(G1), .A3(new_n728), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT99), .Z(new_n956));
  NAND3_X1  g0756(.A1(new_n948), .A2(new_n952), .A3(new_n956), .ZN(G367));
  OAI211_X1 g0757(.A(new_n628), .B(new_n635), .C1(new_n619), .C2(new_n667), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n628), .B2(new_n667), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT108), .ZN(new_n960));
  AND2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n959), .A2(new_n960), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OR2_X1    g0763(.A1(new_n963), .A2(new_n676), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT42), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(KEYINPUT43), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n632), .A2(new_n667), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n649), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n649), .A2(new_n633), .A3(new_n968), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n961), .A2(new_n962), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n549), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n666), .B1(new_n974), .B2(new_n628), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n966), .A2(new_n967), .A3(new_n972), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n972), .A2(new_n967), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n971), .A2(KEYINPUT43), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(new_n965), .C2(new_n975), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n675), .A2(new_n963), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n681), .B(KEYINPUT41), .Z(new_n984));
  NAND2_X1  g0784(.A1(new_n501), .A2(new_n667), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n673), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(new_n676), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(new_n670), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n725), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n973), .A2(new_n678), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT45), .Z(new_n991));
  NOR2_X1   g0791(.A1(new_n973), .A2(new_n678), .ZN(new_n992));
  XNOR2_X1  g0792(.A(KEYINPUT109), .B(KEYINPUT44), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  AOI211_X1 g0794(.A(KEYINPUT110), .B(new_n674), .C1(new_n991), .C2(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(KEYINPUT110), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n675), .A2(new_n996), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n674), .A2(KEYINPUT110), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n991), .A2(new_n997), .A3(new_n994), .A4(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n989), .B1(new_n995), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n984), .B1(new_n1001), .B2(new_n726), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n983), .B1(new_n1002), .B2(new_n731), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n236), .A2(new_n740), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n749), .B1(new_n217), .B2(new_n325), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n732), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n770), .A2(new_n350), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n252), .B1(new_n761), .B2(G317), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n332), .B2(new_n769), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1007), .B(new_n1009), .C1(new_n755), .C2(G311), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT46), .ZN(new_n1011));
  NOR3_X1   g0811(.A1(new_n764), .A2(new_n1011), .A3(new_n485), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1011), .B1(new_n764), .B2(new_n485), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n774), .B2(new_n791), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n1012), .B(new_n1014), .C1(G303), .C2(new_n825), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1010), .B(new_n1015), .C1(new_n787), .C2(new_n782), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n782), .A2(new_n410), .B1(new_n221), .B2(new_n774), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT111), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n252), .B1(new_n770), .B2(new_n251), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT112), .Z(new_n1021));
  INV_X1    g0821(.A(new_n764), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n1022), .A2(G58), .B1(new_n761), .B2(G137), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n768), .A2(G68), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(new_n301), .C2(new_n773), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G143), .B2(new_n755), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1019), .A2(new_n1021), .A3(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n1016), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT47), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1006), .B1(new_n1030), .B2(new_n745), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n972), .A2(new_n748), .ZN(new_n1032));
  AND2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1003), .A2(new_n1034), .ZN(G387));
  INV_X1    g0835(.A(new_n989), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n725), .A2(new_n988), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1036), .A2(new_n681), .A3(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n988), .A2(new_n730), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n732), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n233), .A2(new_n265), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n683), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1041), .A2(new_n739), .B1(new_n1042), .B2(new_n735), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n294), .A2(new_n221), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT50), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n265), .B1(new_n203), .B2(new_n251), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n1045), .A2(new_n1042), .A3(new_n1046), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n1043), .A2(new_n1047), .B1(G107), .B2(new_n217), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1040), .B1(new_n1048), .B2(new_n749), .ZN(new_n1049));
  AOI22_X1  g0849(.A1(G50), .A2(new_n825), .B1(new_n824), .B2(G68), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n363), .B(new_n1007), .C1(G150), .C2(new_n761), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1022), .A2(G77), .ZN(new_n1052));
  OR2_X1    g0852(.A1(new_n769), .A2(new_n325), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1050), .A2(new_n1051), .A3(new_n1052), .A4(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n755), .A2(G159), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT113), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1054), .B(new_n1056), .C1(new_n828), .C2(new_n298), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n770), .A2(new_n485), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n363), .B1(new_n760), .B2(new_n795), .ZN(new_n1059));
  AOI22_X1  g0859(.A1(G303), .A2(new_n824), .B1(new_n825), .B2(G317), .ZN(new_n1060));
  OAI221_X1 g0860(.A(new_n1060), .B1(new_n785), .B2(new_n756), .C1(new_n782), .C2(new_n784), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT48), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n769), .A2(new_n791), .B1(new_n764), .B2(new_n787), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  AOI211_X1 g0866(.A(new_n1058), .B(new_n1059), .C1(new_n1066), .C2(KEYINPUT49), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1066), .A2(KEYINPUT49), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1057), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1049), .B1(new_n1069), .B2(new_n840), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n673), .B2(new_n748), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1039), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1038), .A2(new_n1072), .ZN(G393));
  INV_X1    g0873(.A(new_n995), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1074), .A2(new_n1036), .A3(new_n999), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n681), .A3(new_n1001), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n245), .A2(new_n740), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n749), .B1(new_n350), .B2(new_n217), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n755), .A2(G317), .B1(new_n825), .B2(G311), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT52), .Z(new_n1080));
  OAI221_X1 g0880(.A(new_n363), .B1(new_n760), .B2(new_n785), .C1(new_n332), .C2(new_n770), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n769), .A2(new_n485), .B1(new_n764), .B2(new_n791), .ZN(new_n1082));
  AOI211_X1 g0882(.A(new_n1081), .B(new_n1082), .C1(G294), .C2(new_n824), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n1080), .B(new_n1083), .C1(new_n792), .C2(new_n782), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n755), .A2(G150), .B1(new_n825), .B2(G159), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n1085), .B(KEYINPUT51), .Z(new_n1086));
  OAI22_X1  g0886(.A1(new_n769), .A2(new_n251), .B1(new_n764), .B2(new_n203), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n363), .B1(new_n761), .B2(G143), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1088), .B1(new_n821), .B2(new_n770), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1087), .B(new_n1089), .C1(new_n294), .C2(new_n824), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n1086), .B(new_n1090), .C1(new_n221), .C2(new_n782), .ZN(new_n1091));
  AND2_X1   g0891(.A1(new_n1084), .A2(new_n1091), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n732), .B1(new_n1077), .B2(new_n1078), .C1(new_n1092), .C2(new_n840), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n963), .B2(new_n748), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1074), .A2(new_n999), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1094), .B1(new_n1095), .B2(new_n731), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1076), .A2(new_n1096), .ZN(G390));
  INV_X1    g0897(.A(KEYINPUT117), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n896), .A2(new_n903), .A3(G330), .A4(new_n814), .ZN(new_n1099));
  XNOR2_X1  g0899(.A(new_n1099), .B(KEYINPUT114), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n930), .B1(new_n699), .B2(new_n813), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n927), .B1(new_n1101), .B2(new_n903), .ZN(new_n1102));
  NAND3_X1  g0902(.A1(new_n888), .A2(new_n1102), .A3(new_n895), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n927), .B1(new_n933), .B2(new_n903), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n893), .A2(new_n875), .A3(new_n878), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n925), .B1(new_n1105), .B2(new_n923), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1100), .B(new_n1103), .C1(new_n1104), .C2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT115), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n924), .A2(new_n926), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n940), .B2(new_n927), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1111), .A2(KEYINPUT115), .A3(new_n1103), .A4(new_n1100), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1103), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1099), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n1109), .A2(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n456), .A2(new_n723), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n1116), .B(new_n647), .C1(new_n701), .C2(new_n648), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n903), .B1(new_n723), .B2(new_n814), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n933), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT116), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT116), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n933), .B(new_n1121), .C1(new_n1114), .C2(new_n1118), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1120), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1114), .A2(KEYINPUT114), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1118), .A2(new_n1101), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT114), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1099), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1117), .B1(new_n1123), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(new_n681), .B1(new_n1115), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1109), .A2(new_n1112), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1132));
  AND3_X1   g0932(.A1(new_n1131), .A2(new_n1132), .A3(new_n1129), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1098), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1129), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1131), .A2(new_n1132), .A3(new_n1129), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1137), .A2(KEYINPUT117), .A3(new_n681), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1134), .A2(new_n1139), .ZN(new_n1140));
  INV_X1    g0940(.A(G125), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n252), .B1(new_n760), .B2(new_n1141), .C1(new_n221), .C2(new_n770), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(KEYINPUT54), .B(G143), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n834), .A2(new_n773), .B1(new_n774), .B2(new_n1143), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n1142), .B(new_n1144), .C1(G159), .C2(new_n768), .ZN(new_n1145));
  INV_X1    g0945(.A(KEYINPUT53), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1146), .B1(new_n764), .B2(new_n301), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1022), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1148));
  AOI22_X1  g0948(.A1(new_n755), .A2(G128), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n1145), .B(new_n1149), .C1(new_n782), .C2(new_n831), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n363), .B1(new_n760), .B2(new_n787), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n769), .A2(new_n251), .B1(new_n764), .B2(new_n821), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1151), .B(new_n1152), .C1(G68), .C2(new_n837), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G97), .A2(new_n824), .B1(new_n825), .B2(G116), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1153), .B(new_n1154), .C1(new_n791), .C2(new_n756), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n782), .A2(new_n332), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1150), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n840), .B1(new_n1157), .B2(KEYINPUT118), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(KEYINPUT118), .B2(new_n1157), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1040), .B1(new_n818), .B2(new_n299), .ZN(new_n1160));
  OAI211_X1 g0960(.A(new_n1159), .B(new_n1160), .C1(new_n1106), .C2(new_n747), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1162), .B1(new_n1115), .B2(new_n731), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1140), .A2(new_n1163), .ZN(G378));
  INV_X1    g0964(.A(KEYINPUT57), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n916), .A2(G330), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n911), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n321), .A2(KEYINPUT55), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n320), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n314), .B2(new_n315), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT55), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n307), .A2(new_n863), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT121), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1174), .B(new_n1176), .Z(new_n1177));
  NAND3_X1  g0977(.A1(new_n1169), .A2(new_n1173), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1177), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1180));
  AOI211_X1 g0980(.A(KEYINPUT55), .B(new_n1170), .C1(new_n314), .C2(new_n315), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1179), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1168), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(KEYINPUT104), .B1(new_n941), .B2(new_n928), .ZN(new_n1185));
  AND4_X1   g0985(.A1(KEYINPUT104), .A2(new_n928), .A3(new_n929), .A4(new_n935), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1183), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n911), .A2(new_n1167), .A3(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1184), .A2(new_n1187), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1188), .B1(new_n911), .B2(new_n1167), .ZN(new_n1191));
  AOI211_X1 g0991(.A(new_n1166), .B(new_n1183), .C1(new_n908), .C2(new_n910), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n943), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1117), .B1(new_n1115), .B2(new_n1129), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1165), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1117), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1138), .A2(new_n1197), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1198), .A2(KEYINPUT57), .A3(new_n1190), .A4(new_n1193), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1196), .A2(new_n1199), .A3(new_n681), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1190), .A2(new_n1193), .A3(new_n731), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n732), .B1(new_n819), .B2(G50), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n252), .A2(G41), .ZN(new_n1203));
  AOI211_X1 g1003(.A(G50), .B(new_n1203), .C1(new_n302), .C2(new_n264), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n332), .A2(new_n773), .B1(new_n774), .B2(new_n325), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1024), .B1(new_n202), .B2(new_n770), .C1(new_n791), .C2(new_n760), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n1205), .B(new_n1206), .C1(G116), .C2(new_n755), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1052), .A2(new_n1203), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT119), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1207), .B(new_n1209), .C1(new_n350), .C2(new_n782), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT58), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1204), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n774), .A2(new_n831), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n769), .A2(new_n301), .B1(new_n764), .B2(new_n1143), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(G128), .C2(new_n825), .ZN(new_n1215));
  OAI221_X1 g1015(.A(new_n1215), .B1(new_n1141), .B2(new_n756), .C1(new_n782), .C2(new_n834), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1216), .A2(KEYINPUT59), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n837), .A2(G159), .ZN(new_n1218));
  AOI211_X1 g1018(.A(G33), .B(G41), .C1(new_n761), .C2(G124), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1217), .A2(new_n1218), .A3(new_n1219), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1216), .A2(KEYINPUT59), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1212), .B1(new_n1211), .B2(new_n1210), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1202), .B1(new_n1222), .B2(new_n745), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n1188), .B2(new_n747), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1201), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1200), .A2(new_n1225), .ZN(G375));
  INV_X1    g1026(.A(new_n984), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1122), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n896), .A2(G330), .A3(new_n814), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n939), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1230), .A2(new_n1099), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1121), .B1(new_n1231), .B2(new_n933), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1117), .B(new_n1128), .C1(new_n1228), .C2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1136), .A2(new_n1227), .A3(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n732), .B1(new_n819), .B2(G68), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1053), .B1(new_n350), .B2(new_n764), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n363), .B1(new_n760), .B2(new_n792), .C1(new_n251), .C2(new_n770), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n332), .A2(new_n774), .B1(new_n773), .B2(new_n791), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  OAI221_X1 g1039(.A(new_n1239), .B1(new_n787), .B2(new_n756), .C1(new_n782), .C2(new_n485), .ZN(new_n1240));
  OR2_X1    g1040(.A1(new_n782), .A2(new_n1143), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n756), .A2(new_n834), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n363), .B1(new_n761), .B2(G128), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n202), .B2(new_n770), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n769), .A2(new_n221), .B1(new_n764), .B2(new_n410), .ZN(new_n1245));
  OAI22_X1  g1045(.A1(new_n831), .A2(new_n773), .B1(new_n774), .B2(new_n301), .ZN(new_n1246));
  NOR4_X1   g1046(.A1(new_n1242), .A2(new_n1244), .A3(new_n1245), .A4(new_n1246), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1240), .A2(KEYINPUT122), .B1(new_n1241), .B2(new_n1247), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1248), .B1(KEYINPUT122), .B2(new_n1240), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1235), .B1(new_n1249), .B2(new_n745), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1250), .B(KEYINPUT123), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n746), .B2(new_n939), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1128), .B1(new_n1228), .B2(new_n1232), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1252), .B1(new_n1253), .B2(new_n731), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1234), .A2(new_n1254), .ZN(G381));
  INV_X1    g1055(.A(G387), .ZN(new_n1256));
  INV_X1    g1056(.A(G390), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1038), .A2(new_n802), .A3(new_n1072), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1256), .A2(new_n844), .A3(new_n1257), .A4(new_n1259), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1163), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1261));
  OR4_X1    g1061(.A1(G375), .A2(new_n1260), .A3(G381), .A4(new_n1261), .ZN(G407));
  NAND2_X1  g1062(.A1(new_n1201), .A2(new_n1224), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1198), .A2(new_n1190), .A3(new_n1193), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n682), .B1(new_n1264), .B2(new_n1165), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1263), .B1(new_n1265), .B2(new_n1199), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1261), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n665), .A2(G213), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1267), .A3(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(G407), .A2(G213), .A3(new_n1270), .ZN(G409));
  INV_X1    g1071(.A(KEYINPUT61), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT127), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(G393), .A2(G396), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1273), .B1(new_n1275), .B2(new_n1259), .ZN(new_n1276));
  AND3_X1   g1076(.A1(new_n1003), .A2(new_n1034), .A3(G390), .ZN(new_n1277));
  AOI21_X1  g1077(.A(G390), .B1(new_n1003), .B2(new_n1034), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1276), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G387), .A2(new_n1257), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1003), .A2(new_n1034), .A3(G390), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1274), .A2(KEYINPUT127), .A3(new_n1258), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1276), .A2(new_n1282), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1280), .A2(new_n1281), .A3(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1279), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n682), .B1(new_n1253), .B2(new_n1197), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1123), .A2(KEYINPUT60), .A3(new_n1117), .A4(new_n1128), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT60), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1233), .A2(new_n1288), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1286), .A2(new_n1287), .A3(new_n1289), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(KEYINPUT124), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT124), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1286), .A2(new_n1289), .A3(new_n1292), .A4(new_n1287), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1254), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n844), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1294), .A2(G384), .A3(new_n1254), .ZN(new_n1297));
  OR2_X1    g1097(.A1(new_n1268), .A2(KEYINPUT126), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1269), .A2(G2897), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1299), .A2(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1296), .A2(new_n1297), .A3(new_n1300), .A4(new_n1298), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(G378), .A2(new_n1200), .A3(new_n1225), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1198), .A2(new_n1227), .A3(new_n1190), .A4(new_n1193), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1225), .A2(new_n1306), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n1267), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1269), .B1(new_n1305), .B2(new_n1308), .ZN(new_n1309));
  OAI211_X1 g1109(.A(new_n1272), .B(new_n1285), .C1(new_n1304), .C2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1296), .A2(new_n1297), .ZN(new_n1312));
  AOI211_X1 g1112(.A(new_n1269), .B(new_n1312), .C1(new_n1305), .C2(new_n1308), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(KEYINPUT63), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT125), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1315), .B1(new_n1313), .B2(KEYINPUT63), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1163), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1317), .B1(new_n1134), .B2(new_n1139), .ZN(new_n1318));
  OAI21_X1  g1118(.A(new_n1308), .B1(G375), .B2(new_n1318), .ZN(new_n1319));
  INV_X1    g1119(.A(new_n1312), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1319), .A2(new_n1268), .A3(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT63), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1321), .A2(KEYINPUT125), .A3(new_n1322), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1311), .A2(new_n1314), .A3(new_n1316), .A4(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1321), .A2(KEYINPUT62), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1261), .B1(new_n1225), .B2(new_n1306), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1326), .B1(new_n1266), .B2(G378), .ZN(new_n1327));
  OAI211_X1 g1127(.A(new_n1303), .B(new_n1302), .C1(new_n1327), .C2(new_n1269), .ZN(new_n1328));
  INV_X1    g1128(.A(KEYINPUT62), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1309), .A2(new_n1329), .A3(new_n1320), .ZN(new_n1330));
  NAND4_X1  g1130(.A1(new_n1325), .A2(new_n1328), .A3(new_n1272), .A4(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1285), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1324), .A2(new_n1333), .ZN(G405));
  NAND2_X1  g1134(.A1(G375), .A2(new_n1267), .ZN(new_n1335));
  AND2_X1   g1135(.A1(new_n1335), .A2(new_n1305), .ZN(new_n1336));
  OR2_X1    g1136(.A1(new_n1336), .A2(new_n1312), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1336), .A2(new_n1312), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1337), .A2(new_n1332), .A3(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1332), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1339), .A2(new_n1340), .ZN(G402));
endmodule


