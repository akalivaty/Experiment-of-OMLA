//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT0), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(new_n211), .ZN(new_n218));
  NOR2_X1   g0018(.A1(G58), .A2(G68), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n220), .A2(G50), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(new_n215), .A2(new_n216), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G226), .ZN(new_n225));
  INV_X1    g0025(.A(G77), .ZN(new_n226));
  INV_X1    g0026(.A(G244), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n224), .B1(new_n201), .B2(new_n225), .C1(new_n226), .C2(new_n227), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n213), .B1(new_n228), .B2(new_n231), .ZN(new_n232));
  OAI221_X1 g0032(.A(new_n223), .B1(new_n216), .B2(new_n215), .C1(new_n232), .C2(KEYINPUT1), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT64), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n233), .A2(new_n235), .ZN(G361));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n237), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G232), .ZN(new_n240));
  XOR2_X1   g0040(.A(G250), .B(G257), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT65), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G264), .B(G270), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n240), .B(new_n244), .ZN(G358));
  XNOR2_X1  g0045(.A(G68), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n246), .B(KEYINPUT66), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(G50), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G58), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  AOI22_X1  g0054(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n211), .A2(G33), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n217), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G13), .ZN(new_n262));
  NOR3_X1   g0062(.A1(new_n262), .A2(new_n211), .A3(G1), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(new_n201), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n260), .B1(new_n210), .B2(G20), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n265), .B1(new_n266), .B2(new_n201), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n261), .A2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  OAI21_X1  g0069(.A(KEYINPUT71), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT71), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n261), .A2(new_n271), .A3(new_n267), .A4(KEYINPUT9), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n270), .A2(new_n272), .B1(new_n269), .B2(new_n268), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(G222), .A3(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n280), .A2(KEYINPUT67), .A3(G222), .A4(new_n281), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n281), .B1(new_n278), .B2(new_n279), .ZN(new_n287));
  AND2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n287), .A2(G223), .B1(new_n290), .B2(G77), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n275), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  OAI211_X1 g0092(.A(new_n210), .B(G274), .C1(G41), .C2(G45), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n210), .B1(G41), .B2(G45), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n275), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n293), .B1(new_n295), .B2(new_n225), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G190), .ZN(new_n298));
  OAI21_X1  g0098(.A(G200), .B1(new_n292), .B2(new_n296), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n273), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n273), .A2(new_n298), .A3(new_n302), .A4(new_n299), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n297), .A2(G179), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(new_n297), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(new_n268), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n287), .A2(G238), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n280), .A2(G232), .A3(new_n281), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n290), .A2(G107), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n309), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n293), .B1(new_n295), .B2(new_n227), .ZN(new_n315));
  INV_X1    g0115(.A(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT68), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT68), .ZN(new_n318));
  AOI211_X1 g0118(.A(new_n318), .B(new_n315), .C1(new_n312), .C2(new_n313), .ZN(new_n319));
  NOR2_X1   g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g0120(.A(KEYINPUT70), .B1(new_n320), .B2(G179), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n210), .A2(G20), .ZN(new_n322));
  NAND4_X1  g0122(.A1(new_n322), .A2(new_n259), .A3(G77), .A4(new_n217), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(new_n264), .B2(G77), .ZN(new_n324));
  NAND2_X1  g0124(.A1(G20), .A2(G77), .ZN(new_n325));
  INV_X1    g0125(.A(new_n254), .ZN(new_n326));
  XNOR2_X1  g0126(.A(KEYINPUT15), .B(G87), .ZN(new_n327));
  OAI221_X1 g0127(.A(new_n325), .B1(new_n256), .B2(new_n326), .C1(new_n257), .C2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n324), .B1(new_n328), .B2(new_n260), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(new_n320), .B2(new_n306), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT70), .ZN(new_n331));
  INV_X1    g0131(.A(G179), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n331), .B(new_n332), .C1(new_n317), .C2(new_n319), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n321), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n314), .A2(new_n316), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n318), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n314), .A2(KEYINPUT68), .A3(new_n316), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(G200), .A3(new_n337), .ZN(new_n338));
  OAI21_X1  g0138(.A(G190), .B1(new_n317), .B2(new_n319), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT69), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n329), .B(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  AND4_X1   g0142(.A1(new_n304), .A2(new_n308), .A3(new_n334), .A4(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT17), .ZN(new_n344));
  INV_X1    g0144(.A(new_n260), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n278), .A2(new_n211), .A3(new_n279), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT7), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n211), .A4(new_n279), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n203), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n202), .A2(new_n203), .ZN(new_n351));
  OAI21_X1  g0151(.A(G20), .B1(new_n351), .B2(new_n219), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n254), .A2(G159), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(KEYINPUT16), .B1(new_n350), .B2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT7), .B1(new_n290), .B2(new_n211), .ZN(new_n356));
  INV_X1    g0156(.A(new_n349), .ZN(new_n357));
  OAI21_X1  g0157(.A(G68), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT16), .ZN(new_n359));
  INV_X1    g0159(.A(new_n354), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n345), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n256), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(new_n263), .ZN(new_n364));
  INV_X1    g0164(.A(new_n266), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n364), .B1(new_n365), .B2(new_n363), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g0167(.A(G223), .B(new_n281), .C1(new_n288), .C2(new_n289), .ZN(new_n368));
  OAI211_X1 g0168(.A(G226), .B(G1698), .C1(new_n288), .C2(new_n289), .ZN(new_n369));
  NAND2_X1  g0169(.A1(G33), .A2(G87), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n313), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n275), .A2(G232), .A3(new_n294), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(new_n293), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT75), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(KEYINPUT75), .A3(new_n293), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n372), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(G200), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AND3_X1   g0180(.A1(new_n373), .A2(KEYINPUT75), .A3(new_n293), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT75), .B1(new_n373), .B2(new_n293), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G190), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n383), .A2(new_n384), .A3(new_n372), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n344), .B1(new_n367), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n359), .B1(new_n358), .B2(new_n360), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n350), .A2(KEYINPUT16), .A3(new_n354), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n260), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n366), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n386), .A2(new_n390), .A3(new_n344), .A4(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(KEYINPUT76), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT76), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n367), .A2(new_n394), .A3(new_n344), .A4(new_n386), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n387), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n378), .A2(new_n332), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n306), .B1(new_n383), .B2(new_n372), .ZN(new_n398));
  OAI22_X1  g0198(.A1(new_n362), .A2(new_n366), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  XNOR2_X1  g0199(.A(new_n399), .B(KEYINPUT18), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n396), .A2(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n262), .A2(G1), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(G20), .A3(new_n203), .ZN(new_n403));
  XNOR2_X1  g0203(.A(new_n403), .B(KEYINPUT12), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n203), .B2(new_n365), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n254), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n406), .B1(new_n226), .B2(new_n257), .ZN(new_n407));
  AND3_X1   g0207(.A1(new_n407), .A2(KEYINPUT11), .A3(new_n260), .ZN(new_n408));
  AOI21_X1  g0208(.A(KEYINPUT11), .B1(new_n407), .B2(new_n260), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n405), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n280), .A2(G232), .A3(G1698), .ZN(new_n411));
  OAI211_X1 g0211(.A(G226), .B(new_n281), .C1(new_n288), .C2(new_n289), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G97), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT72), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(KEYINPUT72), .A2(G33), .A3(G97), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n411), .A2(new_n412), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n313), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n295), .A2(KEYINPUT73), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT73), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n421), .B1(new_n275), .B2(new_n294), .ZN(new_n422));
  OAI21_X1  g0222(.A(G238), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n293), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(KEYINPUT13), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT13), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n419), .A2(new_n423), .A3(new_n426), .A4(new_n293), .ZN(new_n427));
  AND3_X1   g0227(.A1(new_n425), .A2(new_n384), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(G200), .B1(new_n425), .B2(new_n427), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n410), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(KEYINPUT74), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT74), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n432), .B(new_n410), .C1(new_n428), .C2(new_n429), .ZN(new_n433));
  INV_X1    g0233(.A(new_n293), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n295), .B(KEYINPUT73), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n434), .B1(new_n435), .B2(G238), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n426), .B1(new_n436), .B2(new_n419), .ZN(new_n437));
  INV_X1    g0237(.A(new_n427), .ZN(new_n438));
  OAI21_X1  g0238(.A(G169), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT14), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT14), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n441), .B(G169), .C1(new_n437), .C2(new_n438), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n425), .A2(G179), .A3(new_n427), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n440), .A2(new_n442), .A3(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n410), .ZN(new_n445));
  AOI22_X1  g0245(.A1(new_n431), .A2(new_n433), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AND3_X1   g0246(.A1(new_n343), .A2(new_n401), .A3(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(G107), .B1(new_n356), .B2(new_n357), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n207), .A2(KEYINPUT6), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT77), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n206), .ZN(new_n451));
  NAND2_X1  g0251(.A1(KEYINPUT77), .A2(G97), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G97), .A2(G107), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT6), .B1(new_n208), .B2(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(G20), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n254), .A2(G77), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n448), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n264), .A2(new_n206), .ZN(new_n459));
  OAI211_X1 g0259(.A(new_n264), .B(new_n345), .C1(G1), .C2(new_n277), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(G97), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n458), .A2(new_n260), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n210), .A2(G45), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(KEYINPUT5), .A2(G41), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G274), .ZN(new_n468));
  INV_X1    g0268(.A(G45), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(G1), .ZN(new_n470));
  INV_X1    g0270(.A(new_n466), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n470), .B1(new_n471), .B2(new_n464), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n275), .ZN(new_n473));
  INV_X1    g0273(.A(G257), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI211_X1 g0275(.A(G244), .B(new_n281), .C1(new_n288), .C2(new_n289), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT78), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT4), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT4), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(G283), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n277), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n483), .B1(new_n287), .B2(G250), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n479), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  AOI211_X1 g0285(.A(G190), .B(new_n475), .C1(new_n485), .C2(new_n313), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n484), .A2(new_n481), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n480), .B1(new_n476), .B2(new_n477), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n313), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n475), .ZN(new_n490));
  AOI21_X1  g0290(.A(G200), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n462), .B1(new_n486), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n458), .A2(new_n260), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n461), .A2(new_n459), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AOI211_X1 g0295(.A(new_n332), .B(new_n475), .C1(new_n485), .C2(new_n313), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n306), .B1(new_n489), .B2(new_n490), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n451), .A2(new_n452), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n499), .A2(new_n211), .A3(G33), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT19), .ZN(new_n501));
  AOI21_X1  g0301(.A(G20), .B1(new_n278), .B2(new_n279), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(G68), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n415), .A2(KEYINPUT19), .A3(new_n416), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT79), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n505), .A3(new_n211), .ZN(new_n506));
  INV_X1    g0306(.A(G87), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n451), .A2(new_n507), .A3(new_n207), .A4(new_n452), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n505), .B1(new_n504), .B2(new_n211), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n260), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n327), .A2(new_n263), .ZN(new_n513));
  OR2_X1    g0313(.A1(new_n460), .A2(new_n327), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n513), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n463), .A2(G250), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n470), .A2(G274), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n313), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g0318(.A(G244), .B(G1698), .C1(new_n288), .C2(new_n289), .ZN(new_n519));
  OAI211_X1 g0319(.A(G238), .B(new_n281), .C1(new_n288), .C2(new_n289), .ZN(new_n520));
  NAND2_X1  g0320(.A1(G33), .A2(G116), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n518), .B1(new_n522), .B2(new_n313), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G179), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n306), .B2(new_n523), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n515), .A2(new_n525), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n511), .A2(new_n260), .B1(new_n263), .B2(new_n327), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n523), .A2(new_n384), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(G200), .B2(new_n523), .ZN(new_n529));
  INV_X1    g0329(.A(new_n460), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(G87), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n527), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  AND4_X1   g0332(.A1(new_n492), .A2(new_n498), .A3(new_n526), .A4(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(KEYINPUT81), .B1(new_n521), .B2(G20), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT81), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n535), .A2(new_n211), .A3(G33), .A4(G116), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT23), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n538), .B1(new_n211), .B2(G107), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND2_X1   g0341(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT22), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n543), .B1(new_n502), .B2(G87), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n211), .B(G87), .C1(new_n288), .C2(new_n289), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(KEYINPUT22), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n542), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT24), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n542), .B(KEYINPUT24), .C1(new_n544), .C2(new_n546), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n549), .A2(new_n260), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n402), .A2(G20), .A3(new_n207), .ZN(new_n552));
  XNOR2_X1  g0352(.A(new_n552), .B(KEYINPUT25), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n553), .B1(new_n530), .B2(G107), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n472), .A2(G264), .A3(new_n275), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT82), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n472), .A2(KEYINPUT82), .A3(G264), .A4(new_n275), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  OAI211_X1 g0359(.A(G250), .B(new_n281), .C1(new_n288), .C2(new_n289), .ZN(new_n560));
  OAI211_X1 g0360(.A(G257), .B(G1698), .C1(new_n288), .C2(new_n289), .ZN(new_n561));
  NAND2_X1  g0361(.A1(G33), .A2(G294), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n313), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n559), .A2(G179), .A3(new_n468), .A4(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n468), .A3(new_n555), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G169), .ZN(new_n567));
  AOI22_X1  g0367(.A1(new_n551), .A2(new_n554), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  AND3_X1   g0368(.A1(new_n564), .A2(new_n468), .A3(new_n555), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n564), .A2(new_n557), .A3(new_n468), .A4(new_n558), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n569), .A2(new_n384), .B1(new_n570), .B2(new_n379), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n550), .A2(new_n260), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n537), .A2(new_n541), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n545), .A2(KEYINPUT22), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n502), .A2(new_n543), .A3(G87), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n573), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n576), .A2(KEYINPUT24), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n554), .B1(new_n572), .B2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(KEYINPUT83), .B1(new_n571), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n570), .A2(new_n379), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n564), .A2(new_n384), .A3(new_n468), .A4(new_n555), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT83), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n551), .A4(new_n554), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n568), .B1(new_n579), .B2(new_n584), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n211), .B1(new_n277), .B2(new_n482), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n451), .A2(new_n452), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(G33), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT80), .ZN(new_n590));
  INV_X1    g0390(.A(G116), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n259), .A2(new_n217), .B1(G20), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n589), .A2(new_n590), .A3(KEYINPUT20), .A4(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(G33), .B1(new_n451), .B2(new_n452), .ZN(new_n594));
  OAI211_X1 g0394(.A(KEYINPUT20), .B(new_n592), .C1(new_n594), .C2(new_n586), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT80), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT20), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n594), .A2(new_n586), .ZN(new_n598));
  INV_X1    g0398(.A(new_n592), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n597), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n593), .A2(new_n596), .A3(new_n600), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n264), .A2(G116), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n602), .B1(new_n530), .B2(G116), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(G264), .B(G1698), .C1(new_n288), .C2(new_n289), .ZN(new_n605));
  OAI211_X1 g0405(.A(G257), .B(new_n281), .C1(new_n288), .C2(new_n289), .ZN(new_n606));
  INV_X1    g0406(.A(G303), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n605), .B(new_n606), .C1(new_n607), .C2(new_n280), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n313), .ZN(new_n609));
  XNOR2_X1  g0409(.A(KEYINPUT5), .B(G41), .ZN(new_n610));
  INV_X1    g0410(.A(new_n217), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n610), .A2(new_n470), .B1(new_n611), .B2(new_n274), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n612), .A2(G270), .B1(G274), .B2(new_n467), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(new_n613), .A3(new_n384), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n609), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n379), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n604), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n306), .B1(new_n609), .B2(new_n613), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT21), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n609), .A2(new_n613), .A3(G179), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n619), .A2(new_n620), .B1(new_n601), .B2(new_n603), .ZN(new_n621));
  AOI21_X1  g0421(.A(KEYINPUT21), .B1(new_n604), .B2(new_n618), .ZN(new_n622));
  NOR3_X1   g0422(.A1(new_n617), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n447), .A2(new_n533), .A3(new_n585), .A4(new_n623), .ZN(G372));
  INV_X1    g0424(.A(new_n334), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n430), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n444), .A2(new_n445), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n396), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OR2_X1    g0428(.A1(new_n628), .A2(new_n400), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n629), .A2(new_n304), .B1(new_n268), .B2(new_n307), .ZN(new_n630));
  INV_X1    g0430(.A(new_n447), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n526), .A2(new_n532), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n632), .B1(new_n633), .B2(new_n498), .ZN(new_n634));
  INV_X1    g0434(.A(new_n498), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n635), .A2(KEYINPUT26), .A3(new_n526), .A4(new_n532), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n492), .A2(new_n498), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n579), .A2(new_n584), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n526), .A2(new_n532), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n604), .A2(new_n618), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT21), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI211_X1 g0443(.A(new_n642), .B(new_n306), .C1(new_n609), .C2(new_n613), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n609), .A2(new_n613), .A3(G179), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n604), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI22_X1  g0446(.A1(new_n569), .A2(new_n306), .B1(new_n570), .B2(new_n332), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n578), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g0448(.A1(new_n643), .A2(new_n646), .A3(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n638), .A2(new_n639), .A3(new_n640), .A4(new_n649), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n637), .A2(new_n650), .A3(new_n526), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n630), .B1(new_n631), .B2(new_n652), .ZN(G369));
  NOR2_X1   g0453(.A1(new_n621), .A2(new_n622), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n402), .ZN(new_n656));
  OR3_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .A3(G20), .ZN(new_n657));
  OAI21_X1  g0457(.A(KEYINPUT27), .B1(new_n656), .B2(G20), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n604), .A2(new_n661), .ZN(new_n662));
  MUX2_X1   g0462(.A(new_n655), .B(new_n623), .S(new_n662), .Z(new_n663));
  XNOR2_X1  g0463(.A(KEYINPUT84), .B(G330), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n578), .A2(new_n661), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n585), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n568), .A2(new_n661), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n666), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n661), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n655), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n568), .A2(new_n673), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n672), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n214), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(new_n210), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n508), .A2(G116), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n682), .A2(new_n683), .B1(new_n222), .B2(new_n681), .ZN(new_n684));
  XOR2_X1   g0484(.A(new_n684), .B(KEYINPUT28), .Z(new_n685));
  INV_X1    g0485(.A(new_n526), .ZN(new_n686));
  AOI22_X1  g0486(.A1(new_n654), .A2(new_n648), .B1(new_n579), .B2(new_n584), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n686), .B1(new_n687), .B2(new_n533), .ZN(new_n688));
  NOR3_X1   g0488(.A1(new_n633), .A2(new_n632), .A3(new_n498), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n689), .B1(KEYINPUT85), .B2(new_n634), .ZN(new_n690));
  AND4_X1   g0490(.A1(KEYINPUT85), .A2(new_n640), .A3(KEYINPUT26), .A4(new_n635), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n688), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n692), .A2(KEYINPUT29), .A3(new_n673), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n651), .A2(new_n673), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT29), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n533), .A2(new_n585), .A3(new_n623), .A4(new_n673), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n564), .A2(new_n557), .A3(new_n558), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n522), .A2(new_n313), .ZN(new_n700));
  INV_X1    g0500(.A(new_n518), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n475), .B1(new_n485), .B2(new_n313), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(new_n645), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT30), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n489), .A2(new_n490), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n523), .A2(G179), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n708), .A2(new_n570), .A3(new_n615), .A4(new_n709), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n703), .A2(new_n704), .A3(KEYINPUT30), .A4(new_n645), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT31), .B1(new_n712), .B2(new_n661), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n698), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(new_n665), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n697), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n685), .B1(new_n719), .B2(G1), .ZN(G364));
  NOR2_X1   g0520(.A1(G13), .A2(G33), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  INV_X1    g0523(.A(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n663), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n217), .B1(G20), .B2(new_n306), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n680), .A2(new_n280), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(G45), .B2(new_n221), .ZN(new_n729));
  XOR2_X1   g0529(.A(new_n729), .B(KEYINPUT88), .Z(new_n730));
  AOI21_X1  g0530(.A(new_n730), .B1(new_n249), .B2(G45), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n214), .A2(new_n280), .ZN(new_n732));
  INV_X1    g0532(.A(G355), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n732), .A2(new_n733), .B1(G116), .B2(new_n214), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n727), .B1(new_n731), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n211), .A2(G13), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT86), .ZN(new_n737));
  AND3_X1   g0537(.A1(new_n737), .A2(KEYINPUT87), .A3(G45), .ZN(new_n738));
  AOI21_X1  g0538(.A(KEYINPUT87), .B1(new_n737), .B2(G45), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n682), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n211), .A2(new_n384), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n744), .A2(new_n379), .A3(G179), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n332), .A2(G200), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(G322), .ZN(new_n749));
  OAI22_X1  g0549(.A1(new_n746), .A2(new_n607), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n211), .A2(G190), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n751), .A2(new_n332), .A3(G200), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n750), .B1(G283), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(G179), .A2(G200), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n755), .A2(G190), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G20), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G294), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n332), .A2(new_n379), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n743), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G326), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n751), .A2(new_n747), .ZN(new_n762));
  INV_X1    g0562(.A(G311), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n760), .A2(new_n761), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n751), .A2(new_n755), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n280), .B(new_n764), .C1(G329), .C2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(KEYINPUT91), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n759), .A2(new_n768), .A3(new_n751), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n768), .B1(new_n759), .B2(new_n751), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(KEYINPUT33), .B(G317), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n754), .A2(new_n758), .A3(new_n767), .A4(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G159), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n765), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT89), .ZN(new_n778));
  OR2_X1    g0578(.A1(new_n778), .A2(KEYINPUT32), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(KEYINPUT32), .ZN(new_n780));
  INV_X1    g0580(.A(new_n757), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(new_n206), .ZN(new_n782));
  OAI22_X1  g0582(.A1(new_n207), .A2(new_n752), .B1(new_n748), .B2(new_n202), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n760), .A2(new_n201), .B1(new_n762), .B2(new_n226), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n779), .A2(new_n780), .A3(new_n785), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n290), .B1(new_n745), .B2(G87), .ZN(new_n787));
  AOI22_X1  g0587(.A1(KEYINPUT90), .A2(new_n787), .B1(new_n772), .B2(G68), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(KEYINPUT90), .B2(new_n787), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n775), .B1(new_n786), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n742), .B1(new_n790), .B2(new_n726), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n735), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n725), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n666), .ZN(new_n794));
  INV_X1    g0594(.A(new_n742), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n663), .A2(new_n665), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n793), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(G396));
  INV_X1    g0600(.A(new_n726), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(new_n722), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n795), .B1(G77), .B2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n748), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n745), .A2(G107), .B1(G294), .B2(new_n805), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n806), .B1(new_n482), .B2(new_n771), .C1(new_n607), .C2(new_n760), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n290), .B1(new_n752), .B2(new_n507), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n762), .A2(new_n591), .B1(new_n765), .B2(new_n763), .ZN(new_n809));
  NOR4_X1   g0609(.A1(new_n807), .A2(new_n782), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n760), .ZN(new_n811));
  INV_X1    g0611(.A(new_n762), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G137), .A2(new_n811), .B1(new_n812), .B2(G159), .ZN(new_n813));
  INV_X1    g0613(.A(G143), .ZN(new_n814));
  INV_X1    g0614(.A(G150), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n813), .B1(new_n814), .B2(new_n748), .C1(new_n815), .C2(new_n771), .ZN(new_n816));
  INV_X1    g0616(.A(KEYINPUT34), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n745), .A2(G50), .B1(G132), .B2(new_n766), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n290), .B1(new_n753), .B2(G68), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n819), .B(new_n820), .C1(new_n202), .C2(new_n781), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n821), .B1(new_n816), .B2(new_n817), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n810), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  OR2_X1    g0623(.A1(new_n673), .A2(new_n329), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n342), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n334), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n321), .A2(new_n330), .A3(new_n333), .A4(new_n673), .ZN(new_n827));
  AND2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n804), .B1(new_n801), .B2(new_n823), .C1(new_n828), .C2(new_n722), .ZN(new_n829));
  INV_X1    g0629(.A(new_n828), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n694), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g0631(.A(new_n831), .B(KEYINPUT92), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n651), .A2(new_n673), .A3(new_n828), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT93), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n651), .A2(new_n828), .A3(KEYINPUT93), .A4(new_n673), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n742), .B1(new_n839), .B2(new_n717), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n838), .A2(new_n718), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n829), .B1(new_n840), .B2(new_n841), .ZN(G384));
  INV_X1    g0642(.A(new_n659), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n843), .B1(new_n362), .B2(new_n366), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n396), .B2(new_n400), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n386), .A2(new_n390), .A3(new_n391), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n847), .A2(new_n399), .A3(new_n844), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT37), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n852), .A2(KEYINPUT97), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n846), .A2(KEYINPUT38), .A3(new_n849), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(KEYINPUT98), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT98), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n846), .A2(new_n856), .A3(KEYINPUT38), .A4(new_n849), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT97), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n850), .A2(new_n858), .A3(new_n851), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n853), .A2(new_n855), .A3(new_n857), .A4(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT39), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n854), .A2(KEYINPUT95), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT95), .ZN(new_n864));
  NAND4_X1  g0664(.A1(new_n846), .A2(new_n864), .A3(KEYINPUT38), .A4(new_n849), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(KEYINPUT96), .B1(new_n850), .B2(new_n851), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT96), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n869), .B(KEYINPUT38), .C1(new_n846), .C2(new_n849), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n867), .A2(new_n871), .A3(KEYINPUT39), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n444), .A2(new_n445), .A3(new_n673), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n862), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n400), .A2(new_n659), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n445), .A2(new_n661), .ZN(new_n877));
  AND2_X1   g0677(.A1(new_n430), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n627), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n446), .B2(new_n877), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n827), .B(KEYINPUT94), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n881), .B1(new_n837), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n867), .A2(new_n871), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n876), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT99), .ZN(new_n887));
  AND3_X1   g0687(.A1(new_n875), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n887), .B1(new_n875), .B2(new_n886), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n693), .A2(new_n447), .A3(new_n696), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT100), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n693), .A2(new_n447), .A3(KEYINPUT100), .A4(new_n696), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n893), .A2(new_n630), .A3(new_n894), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n890), .B(new_n895), .Z(new_n896));
  INV_X1    g0696(.A(KEYINPUT101), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n716), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g0698(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n899), .A2(new_n713), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(KEYINPUT101), .A3(new_n698), .ZN(new_n901));
  NAND4_X1  g0701(.A1(new_n898), .A2(new_n828), .A3(new_n880), .A4(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n860), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(KEYINPUT40), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT102), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(KEYINPUT40), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n902), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n885), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n905), .A2(new_n911), .ZN(new_n912));
  AND4_X1   g0712(.A1(KEYINPUT101), .A2(new_n698), .A3(new_n714), .A4(new_n715), .ZN(new_n913));
  AOI21_X1  g0713(.A(KEYINPUT101), .B1(new_n900), .B2(new_n698), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n447), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n912), .B(new_n916), .Z(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(new_n664), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n896), .A2(new_n918), .B1(new_n210), .B2(new_n737), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n896), .B2(new_n918), .ZN(new_n920));
  OR3_X1    g0720(.A1(new_n221), .A2(new_n226), .A3(new_n351), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n201), .A2(G68), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n210), .B(G13), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n453), .A2(new_n455), .ZN(new_n924));
  OAI211_X1 g0724(.A(G116), .B(new_n218), .C1(new_n924), .C2(KEYINPUT35), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n925), .B1(KEYINPUT35), .B2(new_n924), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n926), .B(KEYINPUT36), .ZN(new_n927));
  OR3_X1    g0727(.A1(new_n920), .A2(new_n923), .A3(new_n927), .ZN(G367));
  NOR2_X1   g0728(.A1(new_n740), .A2(new_n210), .ZN(new_n929));
  INV_X1    g0729(.A(new_n719), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n638), .B1(new_n462), .B2(new_n673), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n635), .A2(new_n661), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n676), .A2(new_n677), .A3(new_n933), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT45), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n934), .B(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n933), .B1(new_n676), .B2(new_n677), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT44), .ZN(new_n938));
  OR2_X1    g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  AOI22_X1  g0739(.A1(new_n672), .A2(KEYINPUT109), .B1(new_n937), .B2(new_n938), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n936), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n672), .A2(KEYINPUT109), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n941), .B(new_n942), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n675), .B(KEYINPUT107), .Z(new_n944));
  NAND2_X1  g0744(.A1(new_n671), .A2(new_n674), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(KEYINPUT108), .B1(new_n946), .B2(new_n666), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT108), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n944), .A2(new_n794), .A3(new_n948), .A4(new_n945), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n946), .A2(new_n666), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n930), .B1(new_n943), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(KEYINPUT106), .B(KEYINPUT41), .Z(new_n955));
  XNOR2_X1  g0755(.A(new_n681), .B(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n929), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n673), .B1(new_n527), .B2(new_n531), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n526), .A2(new_n958), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n959), .B1(new_n640), .B2(new_n958), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT103), .Z(new_n961));
  INV_X1    g0761(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n963));
  OR3_X1    g0763(.A1(new_n937), .A2(KEYINPUT105), .A3(new_n676), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT42), .ZN(new_n965));
  OAI21_X1  g0765(.A(KEYINPUT105), .B1(new_n937), .B2(new_n676), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n635), .B1(new_n492), .B2(new_n568), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n967), .B1(new_n661), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n965), .B1(new_n964), .B2(new_n966), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n963), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n962), .A2(KEYINPUT43), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT104), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n973), .B(new_n963), .C1(new_n969), .C2(new_n970), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n672), .ZN(new_n978));
  INV_X1    g0778(.A(new_n933), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n977), .A2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n975), .A2(new_n980), .A3(new_n976), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n957), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n728), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n244), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n727), .B1(new_n214), .B2(new_n327), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n795), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n746), .A2(new_n591), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(KEYINPUT46), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n207), .B2(new_n781), .ZN(new_n991));
  INV_X1    g0791(.A(G317), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n290), .B1(new_n992), .B2(new_n765), .C1(new_n989), .C2(KEYINPUT46), .ZN(new_n993));
  INV_X1    g0793(.A(G294), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n771), .A2(new_n994), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n499), .A2(new_n753), .B1(new_n812), .B2(G283), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n607), .B2(new_n748), .C1(new_n763), .C2(new_n760), .ZN(new_n997));
  NOR4_X1   g0797(.A1(new_n991), .A2(new_n993), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n280), .B1(new_n746), .B2(new_n202), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n752), .A2(new_n226), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(G143), .B2(new_n811), .ZN(new_n1001));
  INV_X1    g0801(.A(G137), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1001), .B1(new_n201), .B2(new_n762), .C1(new_n1002), .C2(new_n765), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n999), .B(new_n1003), .C1(G159), .C2(new_n772), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n781), .A2(new_n203), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G150), .B2(new_n805), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT110), .Z(new_n1007));
  AOI21_X1  g0807(.A(new_n998), .B1(new_n1004), .B2(new_n1007), .ZN(new_n1008));
  OR2_X1    g0808(.A1(new_n1008), .A2(KEYINPUT47), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n801), .B1(new_n1008), .B2(KEYINPUT47), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n988), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n962), .B2(new_n724), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n984), .A2(new_n1012), .ZN(G387));
  NAND2_X1  g0813(.A1(new_n953), .A2(new_n719), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n952), .A2(new_n930), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1014), .A2(new_n681), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n290), .B1(new_n752), .B2(new_n591), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(G322), .A2(new_n811), .B1(new_n812), .B2(G303), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n992), .B2(new_n748), .C1(new_n771), .C2(new_n763), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  OR2_X1    g0820(.A1(new_n1020), .A2(KEYINPUT48), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1020), .A2(KEYINPUT48), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n745), .A2(G294), .B1(G283), .B2(new_n757), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(KEYINPUT114), .B(KEYINPUT49), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  AOI211_X1 g0826(.A(new_n1017), .B(new_n1026), .C1(G326), .C2(new_n766), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n771), .A2(new_n256), .B1(new_n203), .B2(new_n762), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT113), .ZN(new_n1029));
  XOR2_X1   g0829(.A(KEYINPUT112), .B(G150), .Z(new_n1030));
  AOI22_X1  g0830(.A1(G50), .A2(new_n805), .B1(new_n766), .B2(new_n1030), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(new_n745), .A2(G77), .B1(G97), .B2(new_n753), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n781), .A2(new_n327), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n290), .B(new_n1033), .C1(G159), .C2(new_n811), .ZN(new_n1034));
  AND4_X1   g0834(.A1(new_n1029), .A2(new_n1031), .A3(new_n1032), .A4(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n726), .B1(new_n1027), .B2(new_n1035), .ZN(new_n1036));
  OAI211_X1 g0836(.A(new_n683), .B(new_n469), .C1(new_n203), .C2(new_n226), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT111), .Z(new_n1038));
  NAND2_X1  g0838(.A1(new_n363), .A2(new_n201), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT50), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n728), .B1(new_n1038), .B2(new_n1040), .C1(new_n240), .C2(new_n469), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(G107), .B2(new_n214), .C1(new_n683), .C2(new_n732), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n742), .B1(new_n1042), .B2(new_n727), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1036), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n671), .B2(new_n723), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n929), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1045), .B1(new_n953), .B2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1016), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(KEYINPUT115), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT115), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n1016), .A2(new_n1050), .A3(new_n1047), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1049), .A2(new_n1051), .ZN(G393));
  NOR2_X1   g0852(.A1(new_n952), .A2(new_n930), .ZN(new_n1053));
  OR3_X1    g0853(.A1(new_n1053), .A2(new_n943), .A3(KEYINPUT120), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1053), .A2(new_n943), .ZN(new_n1055));
  AOI21_X1  g0855(.A(KEYINPUT120), .B1(new_n1053), .B2(new_n943), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n1054), .B(new_n681), .C1(new_n1055), .C2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n979), .A2(new_n723), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n727), .B1(new_n214), .B2(new_n588), .C1(new_n985), .C2(new_n252), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n742), .B1(new_n1060), .B2(KEYINPUT116), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(KEYINPUT116), .B2(new_n1060), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n746), .A2(new_n482), .B1(new_n765), .B2(new_n749), .ZN(new_n1063));
  INV_X1    g0863(.A(KEYINPUT117), .ZN(new_n1064));
  OAI221_X1 g0864(.A(new_n290), .B1(new_n207), .B2(new_n752), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n1064), .B2(new_n1063), .ZN(new_n1066));
  XOR2_X1   g0866(.A(new_n1066), .B(KEYINPUT118), .Z(new_n1067));
  OAI22_X1  g0867(.A1(new_n760), .A2(new_n992), .B1(new_n748), .B2(new_n763), .ZN(new_n1068));
  XNOR2_X1  g0868(.A(new_n1068), .B(KEYINPUT52), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n772), .A2(G303), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n812), .A2(G294), .B1(new_n757), .B2(G116), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1067), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n1072), .A2(KEYINPUT119), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n760), .A2(new_n815), .B1(new_n748), .B2(new_n776), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT51), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n772), .A2(G50), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n762), .A2(new_n256), .B1(new_n765), .B2(new_n814), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G68), .B2(new_n745), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n280), .B1(new_n752), .B2(new_n507), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G77), .B2(new_n757), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1072), .A2(KEYINPUT119), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1073), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1062), .B1(new_n1083), .B2(new_n726), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n943), .A2(new_n1046), .B1(new_n1058), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1057), .A2(new_n1085), .ZN(G390));
  AOI21_X1  g0886(.A(new_n882), .B1(new_n835), .B2(new_n836), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n873), .B1(new_n1087), .B2(new_n881), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n855), .A2(new_n857), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n858), .B1(new_n850), .B2(new_n851), .ZN(new_n1090));
  AOI211_X1 g0890(.A(KEYINPUT97), .B(KEYINPUT38), .C1(new_n846), .C2(new_n849), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT39), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1093));
  NOR4_X1   g0893(.A1(new_n866), .A2(new_n868), .A3(new_n870), .A4(new_n861), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1088), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n874), .B1(new_n1089), .B2(new_n1092), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n692), .A2(new_n673), .A3(new_n826), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n827), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n880), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1096), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n880), .A2(new_n665), .A3(new_n716), .A4(new_n828), .ZN(new_n1101));
  AND3_X1   g0901(.A1(new_n1095), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n898), .A2(G330), .A3(new_n828), .A4(new_n901), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1103), .A2(new_n881), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n1095), .B2(new_n1100), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1102), .A2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n915), .A2(G330), .A3(new_n447), .ZN(new_n1107));
  AND4_X1   g0907(.A1(new_n630), .A2(new_n893), .A3(new_n894), .A4(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1087), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n881), .B1(new_n717), .B2(new_n830), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1110), .B1(new_n1103), .B2(new_n881), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n1101), .A2(new_n1097), .A3(new_n827), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1103), .A2(new_n881), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1112), .A2(new_n1115), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1108), .A2(new_n1116), .A3(KEYINPUT121), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT121), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1111), .A2(new_n1109), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n893), .A2(new_n630), .A3(new_n894), .A4(new_n1107), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1118), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1106), .A2(new_n1122), .ZN(new_n1123));
  AND2_X1   g0923(.A1(new_n1117), .A2(new_n1121), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1095), .A2(new_n1100), .A3(new_n1101), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n862), .A2(new_n872), .ZN(new_n1126));
  AOI22_X1  g0926(.A1(new_n1126), .A2(new_n1088), .B1(new_n1099), .B2(new_n1096), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1125), .B1(new_n1127), .B2(new_n1104), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1124), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1123), .A2(new_n1129), .A3(new_n681), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1106), .A2(new_n1046), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n722), .B1(new_n862), .B2(new_n872), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n499), .A2(new_n812), .B1(new_n766), .B2(G294), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1133), .B1(new_n482), .B2(new_n760), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(G107), .B2(new_n772), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n203), .A2(new_n752), .B1(new_n748), .B2(new_n591), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n280), .B(new_n1136), .C1(G87), .C2(new_n745), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(new_n226), .C2(new_n781), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n745), .A2(new_n1030), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT53), .Z(new_n1140));
  OAI221_X1 g0940(.A(new_n280), .B1(new_n752), .B2(new_n201), .C1(new_n781), .C2(new_n776), .ZN(new_n1141));
  INV_X1    g0941(.A(G132), .ZN(new_n1142));
  INV_X1    g0942(.A(G125), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n748), .A2(new_n1142), .B1(new_n765), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(G128), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(KEYINPUT54), .B(G143), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n760), .A2(new_n1145), .B1(new_n762), .B2(new_n1146), .ZN(new_n1147));
  NOR3_X1   g0947(.A1(new_n1141), .A2(new_n1144), .A3(new_n1147), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1140), .B(new_n1148), .C1(new_n1002), .C2(new_n771), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n801), .B1(new_n1138), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n795), .B1(new_n363), .B2(new_n802), .ZN(new_n1151));
  OR3_X1    g0951(.A1(new_n1132), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1130), .A2(new_n1131), .A3(new_n1152), .ZN(G378));
  INV_X1    g0953(.A(new_n681), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1120), .B1(new_n1106), .B2(new_n1122), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n304), .A2(new_n308), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n268), .A2(new_n843), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(new_n1156), .B(new_n1157), .ZN(new_n1158));
  XOR2_X1   g0958(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1159));
  XNOR2_X1  g0959(.A(new_n1158), .B(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1161), .B1(new_n912), .B2(G330), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n915), .A2(new_n828), .A3(new_n880), .A4(new_n908), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n902), .A2(new_n906), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n1163), .A2(new_n1164), .B1(new_n867), .B2(new_n871), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT40), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n860), .B2(new_n903), .ZN(new_n1167));
  OAI211_X1 g0967(.A(G330), .B(new_n1161), .C1(new_n1165), .C2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n1162), .A2(new_n1169), .B1(new_n888), .B2(new_n889), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n875), .A2(new_n886), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(KEYINPUT99), .ZN(new_n1172));
  OAI21_X1  g0972(.A(G330), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n1160), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n875), .A2(new_n886), .A3(new_n887), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1172), .A2(new_n1174), .A3(new_n1175), .A4(new_n1168), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1170), .A2(new_n1176), .ZN(new_n1177));
  OAI21_X1  g0977(.A(KEYINPUT57), .B1(new_n1155), .B2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1108), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT57), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1179), .A2(new_n1180), .A3(new_n1176), .A4(new_n1170), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1154), .B1(new_n1178), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1170), .A2(new_n1176), .A3(new_n1046), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n795), .B1(G50), .B2(new_n802), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G107), .A2(new_n805), .B1(new_n766), .B2(G283), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1185), .B1(new_n327), .B2(new_n762), .C1(new_n771), .C2(new_n206), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n746), .A2(new_n226), .B1(new_n760), .B2(new_n591), .ZN(new_n1187));
  INV_X1    g0987(.A(G41), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1188), .B(new_n290), .C1(new_n752), .C2(new_n202), .ZN(new_n1189));
  NOR4_X1   g0989(.A1(new_n1186), .A2(new_n1005), .A3(new_n1187), .A4(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n290), .A2(new_n1188), .ZN(new_n1191));
  AOI21_X1  g0991(.A(G50), .B1(new_n277), .B2(new_n1188), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n1190), .A2(KEYINPUT58), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G125), .A2(new_n811), .B1(new_n812), .B2(G137), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1194), .B1(new_n815), .B2(new_n781), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1146), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(new_n745), .A2(new_n1196), .B1(G128), .B2(new_n805), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT122), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1195), .B(new_n1198), .C1(G132), .C2(new_n772), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n1200), .A2(KEYINPUT59), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n277), .B(new_n1188), .C1(new_n752), .C2(new_n776), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G124), .B2(new_n766), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT59), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1203), .B1(new_n1199), .B2(new_n1204), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1193), .B1(KEYINPUT58), .B2(new_n1190), .C1(new_n1201), .C2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1184), .B1(new_n1206), .B2(new_n726), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1161), .B2(new_n722), .ZN(new_n1208));
  XOR2_X1   g1008(.A(new_n1208), .B(KEYINPUT123), .Z(new_n1209));
  NAND2_X1  g1009(.A1(new_n1183), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1182), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(G375));
  OAI21_X1  g1012(.A(new_n795), .B1(G68), .B2(new_n802), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n280), .B1(new_n752), .B2(new_n202), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n760), .A2(new_n1142), .B1(new_n748), .B2(new_n1002), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1215), .B(new_n1216), .C1(G50), .C2(new_n757), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(new_n745), .A2(G159), .B1(G128), .B2(new_n766), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1218), .B1(new_n815), .B2(new_n762), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(new_n772), .B2(new_n1196), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n746), .A2(new_n206), .B1(new_n748), .B2(new_n482), .ZN(new_n1221));
  NOR4_X1   g1021(.A1(new_n1221), .A2(new_n1033), .A3(new_n1000), .A4(new_n280), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G107), .A2(new_n812), .B1(new_n766), .B2(G303), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n994), .B2(new_n760), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(G116), .B2(new_n772), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1217), .A2(new_n1220), .B1(new_n1222), .B2(new_n1225), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1214), .B1(new_n801), .B2(new_n1226), .C1(new_n880), .C2(new_n722), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1119), .B2(new_n929), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT124), .Z(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1122), .A2(new_n956), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1229), .B1(new_n1232), .B2(new_n1233), .ZN(G381));
  NOR2_X1   g1034(.A1(G375), .A2(G378), .ZN(new_n1235));
  OR2_X1    g1035(.A1(G387), .A2(G390), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1049), .A2(new_n799), .A3(new_n1051), .ZN(new_n1237));
  NOR4_X1   g1037(.A1(new_n1236), .A2(G384), .A3(G381), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1235), .A2(new_n1238), .ZN(G407));
  INV_X1    g1039(.A(G213), .ZN(new_n1240));
  NOR2_X1   g1040(.A1(new_n1240), .A2(G343), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1235), .A2(new_n1241), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(G407), .A2(new_n1242), .A3(G213), .ZN(G409));
  NAND2_X1  g1043(.A1(G387), .A2(G390), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1236), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(G393), .A2(G396), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(new_n1237), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1245), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1236), .A2(new_n1247), .A3(new_n1244), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1241), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT60), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n681), .B1(new_n1230), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1124), .A2(KEYINPUT60), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1254), .B1(new_n1255), .B2(new_n1231), .ZN(new_n1256));
  INV_X1    g1056(.A(G384), .ZN(new_n1257));
  OR3_X1    g1057(.A1(new_n1256), .A2(new_n1257), .A3(new_n1228), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1257), .B1(new_n1256), .B2(new_n1228), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  AND3_X1   g1060(.A1(new_n1130), .A2(new_n1131), .A3(new_n1152), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1182), .A2(new_n1261), .A3(new_n1210), .ZN(new_n1262));
  NOR3_X1   g1062(.A1(new_n1155), .A2(new_n1177), .A3(new_n956), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1210), .ZN(new_n1265));
  AOI21_X1  g1065(.A(G378), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1252), .B(new_n1260), .C1(new_n1262), .C2(new_n1266), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT126), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1178), .A2(new_n1181), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(new_n681), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1271), .A2(G378), .A3(new_n1265), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1261), .B1(new_n1210), .B2(new_n1263), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1241), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT62), .B1(new_n1274), .B2(new_n1260), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1269), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1252), .B1(new_n1262), .B2(new_n1266), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1241), .A2(G2897), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1258), .A2(new_n1259), .A3(new_n1278), .ZN(new_n1279));
  AOI21_X1  g1079(.A(new_n1278), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT61), .B1(new_n1277), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT126), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1267), .A2(new_n1283), .A3(new_n1268), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1282), .A2(new_n1284), .ZN(new_n1285));
  OAI21_X1  g1085(.A(new_n1251), .B1(new_n1276), .B2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1267), .A2(KEYINPUT125), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(KEYINPUT63), .ZN(new_n1288));
  INV_X1    g1088(.A(new_n1251), .ZN(new_n1289));
  INV_X1    g1089(.A(KEYINPUT63), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1267), .A2(KEYINPUT125), .A3(new_n1290), .ZN(new_n1291));
  NAND4_X1  g1091(.A1(new_n1288), .A2(new_n1289), .A3(new_n1282), .A4(new_n1291), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1286), .A2(new_n1292), .ZN(G405));
  NOR2_X1   g1093(.A1(new_n1262), .A2(KEYINPUT127), .ZN(new_n1294));
  OR2_X1    g1094(.A1(new_n1251), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1251), .A2(new_n1294), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1260), .B1(new_n1211), .B2(G378), .ZN(new_n1297));
  OR3_X1    g1097(.A1(new_n1260), .A2(new_n1211), .A3(G378), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(new_n1295), .A2(new_n1296), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  AND2_X1   g1099(.A1(new_n1251), .A2(new_n1294), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1251), .A2(new_n1294), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1298), .A2(new_n1297), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1300), .A2(new_n1301), .A3(new_n1302), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1299), .A2(new_n1303), .ZN(G402));
endmodule


