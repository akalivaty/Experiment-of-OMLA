//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 1 0 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:13 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n822, new_n823, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202));
  XOR2_X1   g001(.A(G8gat), .B(G36gat), .Z(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT78), .ZN(new_n204));
  XNOR2_X1  g003(.A(G64gat), .B(G92gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  XOR2_X1   g005(.A(KEYINPUT27), .B(G183gat), .Z(new_n207));
  INV_X1    g006(.A(KEYINPUT28), .ZN(new_n208));
  NOR3_X1   g007(.A1(new_n207), .A2(new_n208), .A3(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(G190gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT27), .ZN(new_n211));
  INV_X1    g010(.A(G183gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(KEYINPUT68), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT68), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(G183gat), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n211), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n217));
  OAI211_X1 g016(.A(KEYINPUT70), .B(new_n210), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n218), .A2(new_n208), .ZN(new_n219));
  INV_X1    g018(.A(new_n217), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT68), .B(G183gat), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n220), .B1(new_n221), .B2(new_n211), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(new_n210), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT70), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n209), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(G183gat), .A2(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(KEYINPUT67), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT67), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n230), .A2(G169gat), .A3(G176gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT26), .ZN(new_n234));
  INV_X1    g033(.A(G169gat), .ZN(new_n235));
  INV_X1    g034(.A(G176gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n227), .B1(new_n233), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT71), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI211_X1 g041(.A(KEYINPUT71), .B(new_n227), .C1(new_n233), .C2(new_n239), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT23), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n247), .B1(G169gat), .B2(G176gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT23), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n232), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  AND3_X1   g049(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(G183gat), .A2(G190gat), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT65), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT24), .ZN(new_n255));
  AND3_X1   g054(.A1(new_n227), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n254), .B1(new_n227), .B2(new_n255), .ZN(new_n257));
  OAI21_X1  g056(.A(new_n253), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n250), .B1(new_n258), .B2(KEYINPUT66), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT66), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n253), .B(new_n260), .C1(new_n256), .C2(new_n257), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n246), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n232), .A2(new_n248), .A3(new_n249), .ZN(new_n263));
  AOI21_X1  g062(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n251), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n213), .A2(new_n215), .A3(new_n210), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND4_X1  g066(.A1(new_n263), .A2(KEYINPUT69), .A3(KEYINPUT25), .A4(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT69), .ZN(new_n269));
  AND2_X1   g068(.A1(new_n265), .A2(new_n266), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n232), .A2(KEYINPUT25), .A3(new_n248), .A4(new_n249), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n268), .A2(new_n272), .ZN(new_n273));
  OAI22_X1  g072(.A1(new_n226), .A2(new_n244), .B1(new_n262), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT29), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n274), .A2(new_n275), .B1(G226gat), .B2(G233gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(new_n245), .ZN(new_n278));
  AND2_X1   g077(.A1(new_n268), .A2(new_n272), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n242), .A2(new_n243), .ZN(new_n280));
  INV_X1    g079(.A(new_n209), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n218), .A2(new_n208), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT70), .B1(new_n222), .B2(new_n210), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  AOI22_X1  g083(.A1(new_n278), .A2(new_n279), .B1(new_n280), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(G226gat), .A2(G233gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G197gat), .B(G204gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT22), .ZN(new_n289));
  INV_X1    g088(.A(G211gat), .ZN(new_n290));
  INV_X1    g089(.A(G218gat), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G211gat), .B(G218gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(new_n293), .B(new_n294), .ZN(new_n295));
  NOR3_X1   g094(.A1(new_n276), .A2(new_n287), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n294), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n293), .B(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n286), .B1(new_n285), .B2(KEYINPUT29), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n274), .A2(G226gat), .A3(G233gat), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n298), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(new_n206), .B1(new_n296), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n295), .B1(new_n276), .B2(new_n287), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n299), .A2(new_n298), .A3(new_n300), .ZN(new_n304));
  INV_X1    g103(.A(new_n206), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n302), .A2(KEYINPUT30), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT30), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n303), .A2(new_n304), .A3(new_n308), .A4(new_n305), .ZN(new_n309));
  XNOR2_X1  g108(.A(G1gat), .B(G29gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n310), .B(KEYINPUT0), .ZN(new_n311));
  XNOR2_X1  g110(.A(G57gat), .B(G85gat), .ZN(new_n312));
  XOR2_X1   g111(.A(new_n311), .B(new_n312), .Z(new_n313));
  XOR2_X1   g112(.A(G127gat), .B(G134gat), .Z(new_n314));
  XNOR2_X1  g113(.A(G113gat), .B(G120gat), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n314), .B(KEYINPUT72), .C1(KEYINPUT1), .C2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT72), .ZN(new_n317));
  INV_X1    g116(.A(G113gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G120gat), .ZN(new_n319));
  INV_X1    g118(.A(G120gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G113gat), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT1), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(G127gat), .B(G134gat), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n317), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT73), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n319), .A2(new_n321), .A3(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT1), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n318), .A2(KEYINPUT73), .A3(G120gat), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n326), .A2(new_n327), .A3(new_n328), .A4(new_n323), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n316), .A2(new_n324), .A3(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(G141gat), .A2(G148gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(G141gat), .A2(G148gat), .ZN(new_n332));
  OAI21_X1  g131(.A(KEYINPUT79), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(G141gat), .ZN(new_n334));
  INV_X1    g133(.A(G148gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT79), .ZN(new_n337));
  NAND2_X1  g136(.A1(G141gat), .A2(G148gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT2), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n333), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G155gat), .ZN(new_n342));
  INV_X1    g141(.A(G162gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G155gat), .A2(G162gat), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT80), .B1(new_n331), .B2(new_n332), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT80), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n336), .A2(new_n348), .A3(new_n338), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n345), .B1(new_n344), .B2(KEYINPUT2), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n341), .A2(new_n346), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n330), .A2(KEYINPUT4), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT4), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n341), .A2(new_n346), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n350), .A2(new_n351), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n316), .A2(new_n324), .A3(new_n329), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n354), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT3), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n358), .B1(new_n352), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n357), .A2(KEYINPUT3), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n361), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n357), .A2(KEYINPUT3), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n352), .A2(new_n362), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT81), .A4(new_n358), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n360), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(G225gat), .A2(G233gat), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n369), .A2(KEYINPUT5), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT5), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n330), .A2(new_n352), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n370), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n372), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n377), .B1(new_n369), .B2(new_n370), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n313), .B1(new_n371), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT6), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n365), .A2(new_n368), .ZN(new_n381));
  INV_X1    g180(.A(new_n360), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n381), .A2(new_n370), .A3(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n377), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n313), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n369), .A2(KEYINPUT5), .A3(new_n370), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n379), .A2(new_n380), .A3(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n385), .A2(KEYINPUT6), .A3(new_n387), .A4(new_n386), .ZN(new_n390));
  AOI22_X1  g189(.A1(new_n307), .A2(new_n309), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n295), .B1(new_n364), .B2(KEYINPUT29), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n362), .B1(new_n295), .B2(KEYINPUT29), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n357), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n392), .A2(G228gat), .A3(G233gat), .A4(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G228gat), .A2(G233gat), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n298), .A2(new_n275), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n352), .B1(new_n397), .B2(new_n362), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n298), .B1(new_n367), .B2(new_n275), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G22gat), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n395), .A2(new_n400), .A3(KEYINPUT82), .A4(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G78gat), .B(G106gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT31), .B(G50gat), .ZN(new_n404));
  XOR2_X1   g203(.A(new_n403), .B(new_n404), .Z(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  AND2_X1   g205(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n395), .A2(new_n400), .A3(new_n401), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n401), .B1(new_n395), .B2(new_n400), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n408), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT83), .ZN(new_n412));
  AND3_X1   g211(.A1(new_n407), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n407), .A2(new_n411), .ZN(new_n414));
  INV_X1    g213(.A(new_n409), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n408), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n412), .B1(new_n416), .B2(new_n405), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n413), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n225), .A2(new_n208), .A3(new_n218), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n244), .B1(new_n419), .B2(new_n281), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n262), .A2(new_n273), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n330), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n278), .A2(new_n279), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n280), .A2(new_n284), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n423), .A2(new_n424), .A3(new_n358), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(G227gat), .ZN(new_n427));
  INV_X1    g226(.A(G233gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  XNOR2_X1  g229(.A(KEYINPUT75), .B(KEYINPUT34), .ZN(new_n431));
  AND3_X1   g230(.A1(new_n426), .A2(new_n430), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n431), .B1(new_n426), .B2(new_n430), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n422), .A2(new_n429), .A3(new_n425), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT32), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT74), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n435), .A2(KEYINPUT74), .A3(KEYINPUT32), .ZN(new_n439));
  XNOR2_X1  g238(.A(G15gat), .B(G43gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(G71gat), .B(G99gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(new_n435), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n438), .A2(new_n439), .A3(new_n444), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n435), .B(KEYINPUT32), .C1(new_n443), .C2(new_n442), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n434), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n445), .A2(new_n446), .A3(new_n434), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n391), .A2(new_n418), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT35), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n447), .A2(KEYINPUT76), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n445), .A2(new_n446), .ZN(new_n454));
  INV_X1    g253(.A(new_n434), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n454), .A2(KEYINPUT76), .A3(new_n455), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n453), .A2(new_n456), .A3(new_n449), .A4(new_n418), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n391), .A2(KEYINPUT35), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n452), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n453), .A2(KEYINPUT36), .A3(new_n456), .A4(new_n449), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n448), .A2(new_n449), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT36), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT77), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n445), .A2(new_n446), .A3(new_n434), .ZN(new_n464));
  OAI211_X1 g263(.A(KEYINPUT77), .B(new_n462), .C1(new_n464), .C2(new_n447), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n460), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n417), .A2(new_n414), .ZN(new_n468));
  INV_X1    g267(.A(new_n413), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n307), .A2(new_n388), .A3(new_n309), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT39), .B1(new_n375), .B2(new_n376), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g273(.A(KEYINPUT85), .B(KEYINPUT39), .C1(new_n375), .C2(new_n376), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n474), .B(new_n475), .C1(new_n369), .C2(new_n370), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n381), .A2(new_n382), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT84), .B(KEYINPUT39), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n477), .A2(new_n376), .A3(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n476), .A2(new_n479), .A3(KEYINPUT86), .A4(new_n313), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT87), .ZN(new_n481));
  AND2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  AND3_X1   g281(.A1(new_n476), .A2(new_n313), .A3(new_n479), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT86), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n484), .B1(new_n481), .B2(KEYINPUT40), .ZN(new_n485));
  OAI22_X1  g284(.A1(new_n482), .A2(KEYINPUT40), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n470), .B1(new_n471), .B2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT88), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n303), .A2(new_n304), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT37), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT38), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT37), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n303), .A2(new_n304), .A3(new_n488), .A4(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n490), .A2(new_n491), .A3(new_n493), .A4(new_n206), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT89), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n490), .A2(new_n493), .A3(new_n206), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT38), .ZN(new_n497));
  AND3_X1   g296(.A1(new_n389), .A2(new_n390), .A3(new_n306), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n305), .B1(new_n489), .B2(KEYINPUT37), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT89), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n499), .A2(new_n500), .A3(new_n491), .A4(new_n493), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n495), .A2(new_n497), .A3(new_n498), .A4(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n391), .ZN(new_n503));
  AOI22_X1  g302(.A1(new_n487), .A2(new_n502), .B1(new_n470), .B2(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n459), .B1(new_n467), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G113gat), .B(G141gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(G197gat), .ZN(new_n507));
  XOR2_X1   g306(.A(KEYINPUT11), .B(G169gat), .Z(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XOR2_X1   g308(.A(new_n509), .B(KEYINPUT12), .Z(new_n510));
  INV_X1    g309(.A(KEYINPUT93), .ZN(new_n511));
  XNOR2_X1  g310(.A(G15gat), .B(G22gat), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT16), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n512), .B1(new_n513), .B2(G1gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n514), .B1(G1gat), .B2(new_n512), .ZN(new_n515));
  INV_X1    g314(.A(G8gat), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(G29gat), .A2(G36gat), .ZN(new_n518));
  XNOR2_X1  g317(.A(new_n518), .B(KEYINPUT14), .ZN(new_n519));
  XOR2_X1   g318(.A(KEYINPUT90), .B(G29gat), .Z(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(G36gat), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g320(.A(G43gat), .B(G50gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n522), .A2(KEYINPUT15), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n522), .A2(KEYINPUT15), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n521), .B1(KEYINPUT91), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(KEYINPUT91), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n523), .ZN(new_n528));
  OR3_X1    g327(.A1(new_n526), .A2(KEYINPUT92), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(KEYINPUT92), .B1(new_n526), .B2(new_n528), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n524), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI211_X1 g332(.A(KEYINPUT17), .B(new_n524), .C1(new_n529), .C2(new_n530), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n511), .B(new_n517), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n517), .ZN(new_n536));
  INV_X1    g335(.A(new_n530), .ZN(new_n537));
  NOR3_X1   g336(.A1(new_n526), .A2(KEYINPUT92), .A3(new_n528), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT17), .B1(new_n539), .B2(new_n524), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n531), .A2(new_n532), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n536), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g341(.A(KEYINPUT93), .B1(new_n531), .B2(new_n517), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n535), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(G229gat), .A2(G233gat), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(KEYINPUT18), .A3(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n531), .B(new_n536), .ZN(new_n547));
  XOR2_X1   g346(.A(new_n545), .B(KEYINPUT13), .Z(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  OR2_X1    g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT18), .B1(new_n544), .B2(new_n545), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n510), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT94), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n544), .A2(new_n545), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT18), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(new_n510), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n557), .A2(new_n558), .A3(new_n546), .A4(new_n550), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n553), .A2(new_n554), .A3(new_n559), .ZN(new_n560));
  OAI211_X1 g359(.A(KEYINPUT94), .B(new_n510), .C1(new_n551), .C2(new_n552), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n202), .B1(new_n505), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n456), .A2(new_n449), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n447), .A2(KEYINPUT76), .ZN(new_n565));
  NOR3_X1   g364(.A1(new_n564), .A2(new_n565), .A3(new_n470), .ZN(new_n566));
  INV_X1    g365(.A(new_n458), .ZN(new_n567));
  AOI22_X1  g366(.A1(new_n566), .A2(new_n567), .B1(new_n451), .B2(new_n450), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n564), .A2(new_n565), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n462), .B1(new_n464), .B2(new_n447), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT77), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g371(.A1(KEYINPUT36), .A2(new_n569), .B1(new_n572), .B2(new_n465), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n487), .A2(new_n502), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n503), .A2(new_n470), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n568), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n560), .A2(new_n561), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(KEYINPUT95), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT99), .ZN(new_n581));
  INV_X1    g380(.A(G85gat), .ZN(new_n582));
  INV_X1    g381(.A(G92gat), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND3_X1  g383(.A1(KEYINPUT99), .A2(G85gat), .A3(G92gat), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(KEYINPUT7), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  AOI22_X1  g386(.A1(KEYINPUT8), .A2(new_n587), .B1(new_n582), .B2(new_n583), .ZN(new_n588));
  OAI211_X1 g387(.A(new_n586), .B(new_n588), .C1(KEYINPUT7), .C2(new_n584), .ZN(new_n589));
  XNOR2_X1  g388(.A(G99gat), .B(G106gat), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n589), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n593), .B1(new_n540), .B2(new_n541), .ZN(new_n594));
  XNOR2_X1  g393(.A(G190gat), .B(G218gat), .ZN(new_n595));
  AND2_X1   g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n597), .B1(new_n531), .B2(new_n592), .ZN(new_n598));
  OR3_X1    g397(.A1(new_n594), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n595), .B1(new_n594), .B2(new_n598), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G134gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(new_n343), .ZN(new_n603));
  AND4_X1   g402(.A1(KEYINPUT100), .A2(new_n599), .A3(new_n600), .A4(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT100), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n600), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g405(.A1(new_n606), .A2(new_n603), .B1(new_n599), .B2(new_n600), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(G64gat), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n609), .A2(G57gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(G57gat), .ZN(new_n611));
  INV_X1    g410(.A(G71gat), .ZN(new_n612));
  INV_X1    g411(.A(G78gat), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI22_X1  g413(.A1(new_n610), .A2(new_n611), .B1(new_n614), .B2(KEYINPUT9), .ZN(new_n615));
  XNOR2_X1  g414(.A(G71gat), .B(G78gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(KEYINPUT21), .ZN(new_n618));
  XOR2_X1   g417(.A(G127gat), .B(G155gat), .Z(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(KEYINPUT98), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n618), .B(new_n620), .Z(new_n621));
  AOI21_X1  g420(.A(new_n536), .B1(KEYINPUT21), .B2(new_n617), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(KEYINPUT97), .B(KEYINPUT19), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT20), .ZN(new_n625));
  NAND2_X1  g424(.A1(G231gat), .A2(G233gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n626), .B(KEYINPUT96), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n625), .B(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(G183gat), .B(G211gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n623), .B(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n608), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(G176gat), .B(G204gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n593), .A2(KEYINPUT10), .A3(new_n617), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n589), .A2(new_n591), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n640), .A2(KEYINPUT101), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n617), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n593), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(new_n592), .A3(new_n617), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT10), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI211_X1 g446(.A(KEYINPUT102), .B(KEYINPUT10), .C1(new_n643), .C2(new_n644), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n639), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G230gat), .A2(G233gat), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n650), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n643), .A2(new_n653), .A3(new_n644), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n638), .B1(new_n652), .B2(new_n655), .ZN(new_n656));
  OR2_X1    g455(.A1(new_n655), .A2(KEYINPUT103), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n655), .A2(KEYINPUT103), .ZN(new_n658));
  NAND4_X1  g457(.A1(new_n651), .A2(new_n637), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n634), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g460(.A1(new_n580), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n389), .A2(new_n390), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(G1gat), .ZN(G1324gat));
  INV_X1    g465(.A(new_n662), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n307), .A2(new_n309), .ZN(new_n668));
  XNOR2_X1  g467(.A(KEYINPUT16), .B(G8gat), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n668), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n516), .B1(new_n662), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(KEYINPUT42), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(KEYINPUT42), .B2(new_n670), .ZN(G1325gat));
  OR3_X1    g473(.A1(new_n667), .A2(G15gat), .A3(new_n461), .ZN(new_n675));
  OAI21_X1  g474(.A(G15gat), .B1(new_n667), .B2(new_n467), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(G1326gat));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n470), .ZN(new_n678));
  XNOR2_X1  g477(.A(KEYINPUT43), .B(G22gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  INV_X1    g479(.A(new_n608), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n681), .A2(new_n660), .A3(new_n631), .ZN(new_n682));
  AND2_X1   g481(.A1(new_n580), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n520), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n664), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT45), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n467), .A2(new_n504), .ZN(new_n688));
  AOI211_X1 g487(.A(new_n681), .B(new_n687), .C1(new_n688), .C2(new_n568), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT44), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n577), .A2(new_n608), .B1(KEYINPUT104), .B2(new_n690), .ZN(new_n691));
  OR2_X1    g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n562), .A2(new_n660), .A3(new_n631), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n520), .B1(new_n694), .B2(new_n663), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n686), .A2(new_n695), .ZN(G1328gat));
  INV_X1    g495(.A(G36gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n683), .A2(new_n697), .A3(new_n671), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT46), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G36gat), .B1(new_n694), .B2(new_n668), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n700), .A2(new_n701), .A3(KEYINPUT105), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1329gat));
  NOR2_X1   g505(.A1(new_n461), .A2(G43gat), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n683), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(KEYINPUT107), .ZN(new_n709));
  OAI21_X1  g508(.A(G43gat), .B1(new_n694), .B2(new_n467), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n683), .A2(new_n711), .A3(new_n707), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n709), .A2(new_n710), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT106), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g515(.A(new_n470), .B(new_n693), .C1(new_n689), .C2(new_n691), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G50gat), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n418), .A2(G50gat), .ZN(new_n719));
  AOI211_X1 g518(.A(new_n202), .B(new_n562), .C1(new_n688), .C2(new_n568), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT95), .B1(new_n577), .B2(new_n578), .ZN(new_n721));
  OAI211_X1 g520(.A(new_n682), .B(new_n719), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n718), .A2(KEYINPUT48), .A3(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT108), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n580), .A2(KEYINPUT108), .A3(new_n682), .A4(new_n719), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n718), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT109), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT48), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n728), .B1(new_n727), .B2(new_n729), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n723), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT110), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n734), .B(new_n723), .C1(new_n730), .C2(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(G1331gat));
  INV_X1    g535(.A(new_n660), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n578), .A2(new_n634), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n577), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(new_n663), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g540(.A1(new_n739), .A2(new_n668), .ZN(new_n742));
  NOR2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  AND2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n745), .B1(new_n742), .B2(new_n743), .ZN(G1333gat));
  OAI21_X1  g545(.A(G71gat), .B1(new_n739), .B2(new_n467), .ZN(new_n747));
  INV_X1    g546(.A(new_n461), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n612), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(new_n739), .B2(new_n749), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g550(.A1(new_n739), .A2(new_n418), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(new_n613), .ZN(G1335gat));
  NOR2_X1   g552(.A1(new_n578), .A2(new_n631), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n660), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT111), .ZN(new_n756));
  AND2_X1   g555(.A1(new_n692), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G85gat), .B1(new_n758), .B2(new_n663), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n577), .A2(new_n754), .A3(new_n608), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT51), .Z(new_n761));
  NAND4_X1  g560(.A1(new_n761), .A2(new_n582), .A3(new_n664), .A4(new_n660), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(G1336gat));
  OAI21_X1  g562(.A(G92gat), .B1(new_n758), .B2(new_n668), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n761), .A2(new_n583), .A3(new_n671), .A4(new_n660), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT52), .ZN(G1337gat));
  XNOR2_X1  g566(.A(KEYINPUT112), .B(G99gat), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n761), .A2(new_n748), .A3(new_n660), .A4(new_n768), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n758), .A2(new_n467), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n770), .B2(new_n768), .ZN(G1338gat));
  INV_X1    g570(.A(KEYINPUT53), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n737), .A2(G106gat), .A3(new_n418), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n761), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n692), .A2(new_n756), .A3(new_n470), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT114), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G106gat), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n775), .A2(KEYINPUT114), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n772), .B(new_n774), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n775), .A2(G106gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n774), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n781), .A2(KEYINPUT113), .A3(KEYINPUT53), .ZN(new_n782));
  AOI21_X1  g581(.A(KEYINPUT113), .B1(new_n781), .B2(KEYINPUT53), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(G1339gat));
  INV_X1    g583(.A(new_n659), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n651), .A2(KEYINPUT54), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n653), .B(new_n639), .C1(new_n647), .C2(new_n648), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n651), .A2(KEYINPUT54), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n786), .A2(new_n638), .A3(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT55), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n785), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n786), .A2(KEYINPUT55), .A3(new_n638), .A4(new_n788), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n560), .A2(new_n791), .A3(new_n561), .A4(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n547), .A2(new_n549), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n794), .B1(new_n544), .B2(new_n545), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n509), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n660), .A2(new_n559), .A3(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n608), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n791), .A2(new_n608), .A3(new_n792), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n559), .A2(KEYINPUT116), .A3(new_n796), .ZN(new_n800));
  AOI21_X1  g599(.A(KEYINPUT116), .B1(new_n559), .B2(new_n796), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n799), .A2(new_n800), .A3(new_n801), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n632), .B1(new_n798), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n562), .A2(new_n737), .A3(new_n633), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT115), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n562), .A2(KEYINPUT115), .A3(new_n737), .A4(new_n633), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n663), .B1(new_n803), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n461), .A2(new_n470), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n668), .A3(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(G113gat), .B1(new_n811), .B2(new_n562), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n809), .A2(new_n566), .ZN(new_n813));
  XOR2_X1   g612(.A(new_n813), .B(KEYINPUT117), .Z(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n668), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n562), .A2(G113gat), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT118), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n812), .B1(new_n815), .B2(new_n817), .ZN(G1340gat));
  NOR3_X1   g617(.A1(new_n811), .A2(new_n320), .A3(new_n737), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n814), .A2(new_n668), .A3(new_n660), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(new_n320), .ZN(G1341gat));
  OAI21_X1  g620(.A(G127gat), .B1(new_n811), .B2(new_n632), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n632), .A2(G127gat), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n815), .B2(new_n823), .ZN(G1342gat));
  INV_X1    g623(.A(G134gat), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n681), .A2(new_n671), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n814), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT56), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n814), .A2(new_n829), .A3(new_n825), .A4(new_n826), .ZN(new_n830));
  OAI21_X1  g629(.A(G134gat), .B1(new_n811), .B2(new_n681), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(G1343gat));
  AOI211_X1 g631(.A(new_n573), .B(new_n418), .C1(new_n809), .C2(KEYINPUT119), .ZN(new_n833));
  OR2_X1    g632(.A1(new_n809), .A2(KEYINPUT119), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(new_n668), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n334), .B1(new_n835), .B2(new_n562), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n573), .A2(new_n663), .A3(new_n671), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n803), .A2(new_n808), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(new_n470), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT57), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n418), .B1(new_n803), .B2(new_n808), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT57), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n838), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(G141gat), .A3(new_n578), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n836), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT58), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n836), .A2(KEYINPUT58), .A3(new_n846), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1344gat));
  NOR2_X1   g650(.A1(new_n737), .A2(G148gat), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n833), .A2(new_n668), .A3(new_n834), .A4(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n335), .A2(KEYINPUT59), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n855), .B1(new_n845), .B2(new_n660), .ZN(new_n856));
  XOR2_X1   g655(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n857));
  NAND2_X1  g656(.A1(new_n803), .A2(new_n804), .ZN(new_n858));
  AOI21_X1  g657(.A(KEYINPUT57), .B1(new_n858), .B2(new_n470), .ZN(new_n859));
  AOI211_X1 g658(.A(new_n841), .B(new_n418), .C1(new_n803), .C2(new_n808), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n660), .B(new_n837), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n857), .B1(new_n861), .B2(G148gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n853), .B1(new_n856), .B2(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(KEYINPUT121), .B(new_n853), .C1(new_n856), .C2(new_n862), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(G1345gat));
  NOR3_X1   g666(.A1(new_n835), .A2(G155gat), .A3(new_n632), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n342), .B1(new_n845), .B2(new_n631), .ZN(new_n869));
  OR2_X1    g668(.A1(new_n868), .A2(new_n869), .ZN(G1346gat));
  NAND2_X1  g669(.A1(new_n845), .A2(new_n608), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(G162gat), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n833), .A2(new_n343), .A3(new_n826), .A4(new_n834), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n872), .A2(KEYINPUT122), .A3(new_n873), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1347gat));
  NOR2_X1   g677(.A1(new_n664), .A2(new_n668), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n839), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n810), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n882), .A2(G169gat), .A3(new_n578), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n566), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n235), .B1(new_n884), .B2(new_n562), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n883), .A2(new_n885), .ZN(G1348gat));
  NOR3_X1   g685(.A1(new_n881), .A2(new_n236), .A3(new_n737), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n236), .B1(new_n884), .B2(new_n737), .ZN(new_n888));
  OR2_X1    g687(.A1(new_n888), .A2(KEYINPUT123), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(KEYINPUT123), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(G1349gat));
  AOI21_X1  g690(.A(new_n221), .B1(new_n882), .B2(new_n631), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n884), .A2(new_n207), .A3(new_n632), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT60), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n894), .B(new_n895), .ZN(G1350gat));
  NOR3_X1   g695(.A1(new_n884), .A2(G190gat), .A3(new_n681), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT124), .ZN(new_n898));
  OAI21_X1  g697(.A(G190gat), .B1(new_n881), .B2(new_n681), .ZN(new_n899));
  AND2_X1   g698(.A1(new_n899), .A2(KEYINPUT61), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(KEYINPUT61), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(G1351gat));
  NAND2_X1  g701(.A1(new_n467), .A2(new_n879), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n840), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(G197gat), .B1(new_n904), .B2(new_n578), .ZN(new_n905));
  INV_X1    g704(.A(new_n859), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n903), .B1(new_n906), .B2(new_n844), .ZN(new_n907));
  AND2_X1   g706(.A1(new_n578), .A2(G197gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(G1352gat));
  INV_X1    g708(.A(G204gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n904), .A2(new_n910), .A3(new_n660), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT62), .Z(new_n912));
  INV_X1    g711(.A(new_n903), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n660), .B(new_n913), .C1(new_n859), .C2(new_n860), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n912), .B1(new_n910), .B2(new_n915), .ZN(G1353gat));
  NAND3_X1  g715(.A1(new_n907), .A2(KEYINPUT126), .A3(new_n631), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT126), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n913), .B1(new_n859), .B2(new_n860), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n918), .B1(new_n919), .B2(new_n632), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n917), .A2(G211gat), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(KEYINPUT63), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT63), .ZN(new_n923));
  NAND4_X1  g722(.A1(new_n917), .A2(new_n923), .A3(G211gat), .A4(new_n920), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n904), .A2(new_n290), .A3(new_n631), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n925), .B(KEYINPUT125), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n922), .A2(new_n924), .A3(new_n926), .ZN(G1354gat));
  AOI21_X1  g726(.A(G218gat), .B1(new_n904), .B2(new_n608), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n608), .A2(G218gat), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT127), .Z(new_n930));
  AOI21_X1  g729(.A(new_n928), .B1(new_n907), .B2(new_n930), .ZN(G1355gat));
endmodule


