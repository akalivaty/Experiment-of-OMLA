//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n565, new_n566, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n627, new_n630, new_n632, new_n633,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1233,
    new_n1234, new_n1235;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT64), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI211_X1 g036(.A(G137), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT67), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT3), .B(G2104), .ZN(new_n465));
  NAND4_X1  g040(.A1(new_n465), .A2(KEYINPUT67), .A3(G137), .A4(new_n459), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n459), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n468), .B(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G101), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT66), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OR2_X1    g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(G2105), .B1(new_n473), .B2(new_n477), .ZN(new_n478));
  AND3_X1   g053(.A1(new_n467), .A2(new_n471), .A3(new_n478), .ZN(G160));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  AOI21_X1  g057(.A(G2105), .B1(new_n475), .B2(new_n476), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  XNOR2_X1  g059(.A(new_n484), .B(KEYINPUT69), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n459), .B1(new_n475), .B2(new_n476), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n482), .B(new_n485), .C1(G124), .C2(new_n486), .ZN(G162));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT70), .ZN(new_n490));
  OAI21_X1  g065(.A(G2105), .B1(new_n490), .B2(G114), .ZN(new_n491));
  INV_X1    g066(.A(G114), .ZN(new_n492));
  NOR2_X1   g067(.A1(new_n492), .A2(KEYINPUT70), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n489), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  OAI211_X1 g071(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT4), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n465), .A2(new_n499), .A3(G138), .A4(new_n459), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n496), .B1(new_n498), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G62), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n502), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n508));
  INV_X1    g083(.A(G75), .ZN(new_n509));
  OAI22_X1  g084(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n504), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n505), .A2(new_n506), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n511), .A2(new_n508), .A3(G62), .ZN(new_n512));
  INV_X1    g087(.A(new_n512), .ZN(new_n513));
  OAI21_X1  g088(.A(G651), .B1(new_n510), .B2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT6), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n517), .A2(KEYINPUT71), .ZN(new_n518));
  OAI21_X1  g093(.A(G651), .B1(new_n516), .B2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n505), .A2(new_n506), .B1(KEYINPUT6), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n519), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n517), .A2(KEYINPUT71), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n520), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n520), .A2(KEYINPUT6), .ZN(new_n527));
  AND2_X1   g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT5), .A2(G543), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(KEYINPUT72), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g106(.A(KEYINPUT73), .B(G88), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n523), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g108(.A(G543), .B1(new_n517), .B2(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n524), .A2(new_n525), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n534), .B1(new_n535), .B2(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G50), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n514), .A2(new_n533), .A3(new_n537), .ZN(G303));
  INV_X1    g113(.A(G303), .ZN(G166));
  NAND3_X1  g114(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n540));
  XOR2_X1   g115(.A(new_n540), .B(KEYINPUT7), .Z(new_n541));
  AND3_X1   g116(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n542));
  AOI211_X1 g117(.A(new_n541), .B(new_n542), .C1(G51), .C2(new_n536), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n523), .A2(new_n531), .A3(G89), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND2_X1  g121(.A1(G77), .A2(G543), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n528), .A2(new_n529), .ZN(new_n548));
  INV_X1    g123(.A(G64), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI22_X1  g125(.A1(G651), .A2(new_n550), .B1(new_n536), .B2(G52), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n523), .A2(new_n531), .A3(G90), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(G301));
  INV_X1    g128(.A(G301), .ZN(G171));
  AOI22_X1  g129(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(new_n520), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n523), .A2(new_n531), .A3(G81), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n536), .A2(G43), .ZN(new_n558));
  AND3_X1   g133(.A1(new_n557), .A2(KEYINPUT75), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g134(.A(KEYINPUT75), .B1(new_n557), .B2(new_n558), .ZN(new_n560));
  OAI21_X1  g135(.A(new_n556), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G860), .ZN(G153));
  NAND4_X1  g138(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT8), .ZN(new_n566));
  NAND4_X1  g141(.A1(G319), .A2(G483), .A3(G661), .A4(new_n566), .ZN(G188));
  INV_X1    g142(.A(new_n534), .ZN(new_n568));
  XNOR2_X1  g143(.A(KEYINPUT71), .B(KEYINPUT6), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n568), .B(G53), .C1(new_n569), .C2(new_n520), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT9), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n573));
  AOI21_X1  g148(.A(new_n573), .B1(new_n505), .B2(new_n506), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n548), .A2(new_n573), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n572), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  AND2_X1   g152(.A1(G78), .A2(G543), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n523), .A2(new_n531), .A3(G91), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n571), .A2(new_n579), .A3(new_n580), .ZN(G299));
  NAND2_X1  g156(.A1(new_n536), .A2(G49), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n511), .B2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n523), .A2(new_n531), .A3(G87), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT77), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n523), .A2(new_n531), .A3(new_n587), .A4(G87), .ZN(new_n588));
  AOI21_X1  g163(.A(new_n584), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G288));
  NAND3_X1  g165(.A1(new_n523), .A2(new_n531), .A3(G86), .ZN(new_n591));
  OAI21_X1  g166(.A(G61), .B1(new_n528), .B2(new_n529), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(G48), .A2(new_n536), .B1(new_n594), .B2(G651), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(G305));
  NAND2_X1  g171(.A1(G72), .A2(G543), .ZN(new_n597));
  INV_X1    g172(.A(G60), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n548), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n599), .A2(G651), .ZN(new_n600));
  XOR2_X1   g175(.A(KEYINPUT78), .B(G85), .Z(new_n601));
  NAND3_X1  g176(.A1(new_n523), .A2(new_n531), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n536), .A2(G47), .ZN(new_n603));
  AND2_X1   g178(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n604), .A2(KEYINPUT79), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n604), .A2(KEYINPUT79), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(new_n606), .B2(new_n607), .ZN(G290));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NOR2_X1   g184(.A1(G301), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n523), .A2(new_n531), .A3(G92), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g188(.A1(new_n523), .A2(new_n531), .A3(KEYINPUT10), .A4(G92), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n511), .A2(KEYINPUT76), .ZN(new_n616));
  OAI21_X1  g191(.A(G66), .B1(new_n616), .B2(new_n574), .ZN(new_n617));
  NAND2_X1  g192(.A1(G79), .A2(G543), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  AOI22_X1  g194(.A1(new_n619), .A2(G651), .B1(G54), .B2(new_n536), .ZN(new_n620));
  AND3_X1   g195(.A1(new_n615), .A2(new_n620), .A3(KEYINPUT80), .ZN(new_n621));
  AOI21_X1  g196(.A(KEYINPUT80), .B1(new_n615), .B2(new_n620), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g198(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n610), .B1(new_n624), .B2(new_n609), .ZN(G284));
  AOI21_X1  g200(.A(new_n610), .B1(new_n624), .B2(new_n609), .ZN(G321));
  NAND2_X1  g201(.A1(G299), .A2(new_n609), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n627), .B1(G168), .B2(new_n609), .ZN(G297));
  OAI21_X1  g203(.A(new_n627), .B1(G168), .B2(new_n609), .ZN(G280));
  NOR2_X1   g204(.A1(new_n623), .A2(G559), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n630), .B1(G860), .B2(new_n624), .ZN(G148));
  NAND2_X1  g206(.A1(new_n561), .A2(new_n609), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n632), .B1(new_n630), .B2(new_n609), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT81), .ZN(G323));
  XNOR2_X1  g209(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g210(.A1(new_n470), .A2(new_n465), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(new_n638), .B(KEYINPUT13), .Z(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g215(.A1(new_n640), .A2(G2100), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT82), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n483), .A2(G135), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n486), .A2(G123), .ZN(new_n644));
  OR2_X1    g219(.A1(G99), .A2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n645), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(G2096), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n648), .B1(new_n640), .B2(G2100), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n642), .A2(new_n649), .ZN(G156));
  INV_X1    g225(.A(KEYINPUT84), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2427), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2430), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT83), .ZN(new_n658));
  INV_X1    g233(.A(G1341), .ZN(new_n659));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n660));
  NAND4_X1  g235(.A1(new_n655), .A2(new_n660), .A3(KEYINPUT14), .A4(new_n656), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n658), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n659), .B1(new_n658), .B2(new_n661), .ZN(new_n664));
  OAI21_X1  g239(.A(G1348), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n664), .ZN(new_n666));
  INV_X1    g241(.A(G1348), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n666), .A2(new_n667), .A3(new_n662), .ZN(new_n668));
  XOR2_X1   g243(.A(G2451), .B(G2454), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT16), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2443), .B(G2446), .ZN(new_n671));
  XOR2_X1   g246(.A(new_n670), .B(new_n671), .Z(new_n672));
  NAND3_X1  g247(.A1(new_n665), .A2(new_n668), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n673), .A2(G14), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n672), .B1(new_n665), .B2(new_n668), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n651), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n675), .ZN(new_n677));
  NAND4_X1  g252(.A1(new_n677), .A2(KEYINPUT84), .A3(G14), .A4(new_n673), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n676), .A2(new_n678), .ZN(G401));
  INV_X1    g254(.A(KEYINPUT18), .ZN(new_n680));
  XOR2_X1   g255(.A(G2084), .B(G2090), .Z(new_n681));
  XNOR2_X1  g256(.A(G2067), .B(G2678), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(KEYINPUT17), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n681), .A2(new_n682), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n680), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XOR2_X1   g261(.A(KEYINPUT85), .B(G2100), .Z(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(G2072), .B(G2078), .Z(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n683), .B2(KEYINPUT18), .ZN(new_n690));
  XOR2_X1   g265(.A(new_n690), .B(G2096), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n688), .B(new_n691), .ZN(G227));
  XOR2_X1   g267(.A(G1971), .B(G1976), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT19), .ZN(new_n694));
  XOR2_X1   g269(.A(G1956), .B(G2474), .Z(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  AND2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(KEYINPUT86), .B(KEYINPUT20), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n695), .A2(new_n696), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n697), .A2(new_n701), .ZN(new_n702));
  MUX2_X1   g277(.A(new_n702), .B(new_n701), .S(new_n694), .Z(new_n703));
  NOR2_X1   g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(G1991), .B(G1996), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  XOR2_X1   g282(.A(G1981), .B(G1986), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT87), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n707), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(G229));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G24), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n604), .A2(KEYINPUT79), .ZN(new_n716));
  AOI22_X1  g291(.A1(new_n716), .A2(new_n605), .B1(G651), .B2(new_n599), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n715), .B1(new_n717), .B2(new_n714), .ZN(new_n718));
  INV_X1    g293(.A(G1986), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n720), .A2(KEYINPUT88), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n714), .A2(G23), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n589), .B2(new_n714), .ZN(new_n723));
  XNOR2_X1  g298(.A(KEYINPUT33), .B(G1976), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n714), .A2(G22), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G166), .B2(new_n714), .ZN(new_n727));
  INV_X1    g302(.A(G1971), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G6), .B(G305), .S(G16), .Z(new_n730));
  XOR2_X1   g305(.A(KEYINPUT32), .B(G1981), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n725), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT89), .B(KEYINPUT34), .Z(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G29), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G25), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n483), .A2(G131), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n486), .A2(G119), .ZN(new_n739));
  OR2_X1    g314(.A1(G95), .A2(G2105), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n740), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n737), .B1(new_n743), .B2(new_n736), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT35), .B(G1991), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n720), .A2(KEYINPUT88), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n721), .A2(new_n735), .A3(new_n746), .A4(new_n747), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT36), .Z(new_n749));
  NOR2_X1   g324(.A1(G29), .A2(G35), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G162), .B2(G29), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT29), .Z(new_n752));
  INV_X1    g327(.A(G2090), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n714), .A2(G20), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(G299), .B2(G16), .ZN(new_n758));
  INV_X1    g333(.A(G1956), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT24), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n736), .B1(new_n761), .B2(G34), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(KEYINPUT96), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n762), .A2(KEYINPUT96), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n761), .B2(G34), .ZN(new_n765));
  AOI22_X1  g340(.A1(G160), .A2(G29), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT97), .ZN(new_n767));
  INV_X1    g342(.A(G2084), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n754), .A2(new_n760), .A3(new_n769), .ZN(new_n770));
  OAI22_X1  g345(.A1(new_n752), .A2(new_n753), .B1(new_n759), .B2(new_n758), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n736), .A2(G26), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT28), .Z(new_n773));
  NAND2_X1  g348(.A1(new_n486), .A2(G128), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT94), .ZN(new_n775));
  OAI21_X1  g350(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n776));
  INV_X1    g351(.A(G116), .ZN(new_n777));
  AOI21_X1  g352(.A(new_n776), .B1(new_n777), .B2(G2105), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n778), .B1(new_n483), .B2(G140), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n773), .B1(new_n780), .B2(G29), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2067), .ZN(new_n782));
  NOR2_X1   g357(.A1(G5), .A2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT99), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G301), .B2(new_n714), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G1961), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n714), .A2(G21), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(G168), .B2(new_n714), .ZN(new_n788));
  OAI211_X1 g363(.A(new_n782), .B(new_n786), .C1(G1966), .C2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n736), .A2(G33), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT95), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT25), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n483), .A2(G139), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n465), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n459), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n790), .B1(new_n797), .B2(new_n736), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n798), .B(G2072), .Z(new_n799));
  NAND2_X1  g374(.A1(new_n736), .A2(G27), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G164), .B2(new_n736), .ZN(new_n801));
  INV_X1    g376(.A(G2078), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n788), .A2(G1966), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n736), .A2(G32), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n470), .A2(G105), .B1(G141), .B2(new_n483), .ZN(new_n806));
  NAND3_X1  g381(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT26), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G129), .B2(new_n486), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n805), .B1(new_n811), .B2(new_n736), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT27), .B(G1996), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT31), .B(G11), .ZN(new_n815));
  XOR2_X1   g390(.A(KEYINPUT30), .B(G28), .Z(new_n816));
  OAI21_X1  g391(.A(new_n815), .B1(new_n816), .B2(G29), .ZN(new_n817));
  OR2_X1    g392(.A1(new_n647), .A2(new_n736), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(KEYINPUT98), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(KEYINPUT98), .B2(new_n818), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n799), .A2(new_n803), .A3(new_n804), .A4(new_n821), .ZN(new_n822));
  NOR4_X1   g397(.A1(new_n770), .A2(new_n771), .A3(new_n789), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(G4), .A2(G16), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n624), .B2(G16), .ZN(new_n825));
  XOR2_X1   g400(.A(KEYINPUT90), .B(G1348), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT91), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n825), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n714), .A2(G19), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT92), .Z(new_n830));
  OAI21_X1  g405(.A(new_n830), .B1(new_n562), .B2(new_n714), .ZN(new_n831));
  XOR2_X1   g406(.A(KEYINPUT93), .B(G1341), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n831), .B(new_n832), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n823), .A2(new_n828), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n749), .A2(new_n834), .ZN(G311));
  OR2_X1    g410(.A1(new_n749), .A2(new_n834), .ZN(G150));
  NAND2_X1  g411(.A1(new_n624), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  NAND2_X1  g413(.A1(G80), .A2(G543), .ZN(new_n839));
  INV_X1    g414(.A(G67), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n548), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g416(.A1(G651), .A2(new_n841), .B1(new_n536), .B2(G55), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n523), .A2(new_n531), .A3(G93), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n561), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(new_n844), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n846), .B(new_n556), .C1(new_n559), .C2(new_n560), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n838), .B(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT39), .ZN(new_n850));
  AOI21_X1  g425(.A(G860), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n851), .B1(new_n850), .B2(new_n849), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n844), .A2(G860), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n853), .B(KEYINPUT37), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n852), .A2(new_n854), .ZN(G145));
  NAND2_X1  g430(.A1(new_n483), .A2(G142), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n486), .A2(G130), .ZN(new_n857));
  OR2_X1    g432(.A1(G106), .A2(G2105), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n858), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n638), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n638), .A2(new_n860), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n742), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n638), .A2(new_n860), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n865), .A2(new_n743), .A3(new_n861), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT102), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n864), .A2(KEYINPUT102), .A3(new_n866), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n780), .A2(new_n810), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n780), .A2(new_n810), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n797), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n874), .ZN(new_n876));
  INV_X1    g451(.A(new_n797), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n876), .A2(new_n877), .A3(new_n872), .ZN(new_n878));
  XNOR2_X1  g453(.A(G164), .B(KEYINPUT101), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n875), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n875), .A2(new_n878), .ZN(new_n881));
  INV_X1    g456(.A(new_n879), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n871), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n880), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n879), .B1(new_n875), .B2(new_n878), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n870), .B(new_n869), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(G160), .B(new_n647), .ZN(new_n889));
  XNOR2_X1  g464(.A(G162), .B(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(G37), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n883), .A2(new_n880), .ZN(new_n893));
  INV_X1    g468(.A(new_n867), .ZN(new_n894));
  AOI21_X1  g469(.A(KEYINPUT103), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n896));
  AOI211_X1 g471(.A(new_n896), .B(new_n867), .C1(new_n883), .C2(new_n880), .ZN(new_n897));
  OAI211_X1 g472(.A(new_n884), .B(new_n892), .C1(new_n895), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n891), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g475(.A1(new_n717), .A2(G288), .ZN(new_n901));
  NAND2_X1  g476(.A1(G290), .A2(new_n589), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(G303), .B(G305), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT42), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT42), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n906), .A2(new_n910), .A3(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n630), .B(new_n848), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n615), .A2(new_n620), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n571), .A2(new_n579), .A3(new_n580), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT104), .ZN(new_n919));
  NAND3_X1  g494(.A1(G299), .A2(new_n615), .A3(new_n620), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND4_X1  g496(.A1(G299), .A2(new_n615), .A3(new_n620), .A4(KEYINPUT104), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n915), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n920), .ZN(new_n924));
  AOI21_X1  g499(.A(G299), .B1(new_n615), .B2(new_n620), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n915), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(KEYINPUT105), .B(new_n915), .C1(new_n924), .C2(new_n925), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n914), .B(KEYINPUT106), .C1(new_n923), .C2(new_n930), .ZN(new_n931));
  OR2_X1    g506(.A1(new_n630), .A2(new_n848), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n630), .A2(new_n848), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n921), .A2(new_n922), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n931), .A2(new_n936), .ZN(new_n937));
  OR2_X1    g512(.A1(new_n930), .A2(new_n923), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT106), .B1(new_n938), .B2(new_n914), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n913), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n938), .A2(new_n914), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n943), .A2(new_n936), .A3(new_n931), .A4(new_n912), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(G868), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n846), .A2(G868), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n609), .B1(new_n940), .B2(new_n944), .ZN(new_n951));
  OAI21_X1  g526(.A(KEYINPUT107), .B1(new_n951), .B2(new_n948), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n952), .ZN(G295));
  NAND2_X1  g528(.A1(new_n946), .A2(new_n949), .ZN(G331));
  NAND2_X1  g529(.A1(new_n557), .A2(new_n558), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT75), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n557), .A2(KEYINPUT75), .A3(new_n558), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n846), .B1(new_n959), .B2(new_n556), .ZN(new_n960));
  INV_X1    g535(.A(new_n847), .ZN(new_n961));
  OAI21_X1  g536(.A(G171), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n845), .A2(G301), .A3(new_n847), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(G168), .A3(new_n963), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n845), .A2(G301), .A3(new_n847), .ZN(new_n965));
  AOI21_X1  g540(.A(G301), .B1(new_n845), .B2(new_n847), .ZN(new_n966));
  OAI21_X1  g541(.A(G286), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n964), .B(new_n967), .C1(new_n930), .C2(new_n923), .ZN(new_n968));
  NOR3_X1   g543(.A1(new_n965), .A2(new_n966), .A3(G286), .ZN(new_n969));
  AOI21_X1  g544(.A(G168), .B1(new_n962), .B2(new_n963), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n935), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(new_n971), .A3(new_n908), .ZN(new_n972));
  INV_X1    g547(.A(G37), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n908), .B1(new_n968), .B2(new_n971), .ZN(new_n975));
  OAI21_X1  g550(.A(KEYINPUT43), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n934), .B1(new_n967), .B2(new_n964), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT108), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n908), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n915), .B1(new_n918), .B2(new_n920), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n934), .B2(new_n915), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n981), .A2(new_n967), .A3(new_n964), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n971), .A2(KEYINPUT108), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n979), .A2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT43), .ZN(new_n985));
  NAND4_X1  g560(.A1(new_n984), .A2(new_n985), .A3(new_n973), .A4(new_n972), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n976), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n985), .B1(new_n974), .B2(new_n975), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n984), .A2(new_n973), .A3(new_n972), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n988), .B1(new_n989), .B2(new_n985), .ZN(new_n990));
  MUX2_X1   g565(.A(new_n987), .B(new_n990), .S(KEYINPUT44), .Z(G397));
  AND4_X1   g566(.A1(G40), .A2(new_n467), .A3(new_n471), .A4(new_n478), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n498), .A2(new_n500), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n490), .A2(G114), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n492), .A2(KEYINPUT70), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n995), .A2(new_n996), .A3(G2105), .ZN(new_n997));
  AOI22_X1  g572(.A1(new_n486), .A2(G126), .B1(new_n997), .B2(new_n489), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(G1384), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n992), .A2(new_n993), .A3(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT109), .ZN(new_n1003));
  OR2_X1    g578(.A1(new_n780), .A2(G2067), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n780), .A2(G2067), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1004), .A2(new_n811), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G1996), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n992), .A2(new_n1001), .A3(new_n993), .A4(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT46), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT47), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n717), .A2(new_n719), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1013), .A2(new_n1002), .ZN(new_n1014));
  XNOR2_X1  g589(.A(new_n1014), .B(KEYINPUT48), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1009), .A2(new_n810), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1004), .B(new_n1005), .C1(new_n1008), .C2(new_n811), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1016), .B1(new_n1003), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n743), .A2(new_n745), .ZN(new_n1019));
  AND2_X1   g594(.A1(new_n743), .A2(new_n745), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1003), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1012), .B1(new_n1015), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(new_n1004), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1023), .B1(new_n1003), .B2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT126), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n467), .A2(new_n471), .A3(new_n478), .A4(G40), .ZN(new_n1028));
  OAI21_X1  g603(.A(G8), .B1(new_n1001), .B2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n520), .B1(new_n592), .B2(new_n593), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n1031));
  OAI21_X1  g606(.A(G1981), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n591), .A2(new_n595), .A3(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1032), .B1(new_n591), .B2(new_n595), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1029), .B1(new_n1035), .B2(KEYINPUT49), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1032), .ZN(new_n1038));
  NAND2_X1  g613(.A1(G305), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n591), .A2(new_n595), .A3(new_n1032), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT49), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1037), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AOI211_X1 g618(.A(KEYINPUT112), .B(KEYINPUT49), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1036), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT110), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1046), .A2(KEYINPUT55), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  NAND3_X1  g623(.A1(G303), .A2(G8), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g624(.A(G8), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT74), .B1(new_n548), .B2(new_n502), .ZN(new_n1051));
  OAI211_X1 g626(.A(new_n1051), .B(new_n512), .C1(new_n509), .C2(new_n504), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1052), .A2(G651), .B1(G50), .B2(new_n536), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1050), .B1(new_n1053), .B2(new_n533), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1049), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1028), .B1(new_n1001), .B2(new_n993), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n999), .A2(KEYINPUT45), .A3(new_n1000), .ZN(new_n1058));
  AOI21_X1  g633(.A(G1971), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1060));
  AOI21_X1  g635(.A(G1384), .B1(new_n994), .B2(new_n998), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT50), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AND4_X1   g638(.A1(new_n753), .A2(new_n1060), .A3(new_n992), .A4(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1056), .B(G8), .C1(new_n1059), .C2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT52), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(new_n589), .B2(G1976), .ZN(new_n1067));
  INV_X1    g642(.A(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1976), .ZN(new_n1069));
  AOI211_X1 g644(.A(new_n1069), .B(new_n584), .C1(new_n586), .C2(new_n588), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(new_n1029), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1068), .A2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT52), .B1(new_n1070), .B2(new_n1029), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1045), .A2(new_n1065), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1062), .B1(new_n999), .B2(new_n1000), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT114), .B1(new_n1075), .B2(new_n1028), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n1077));
  OAI211_X1 g652(.A(new_n992), .B(new_n1077), .C1(new_n1062), .C2(new_n1061), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1076), .A2(new_n1078), .A3(new_n753), .A4(new_n1063), .ZN(new_n1079));
  OAI21_X1  g654(.A(new_n993), .B1(G164), .B2(G1384), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(new_n992), .A3(new_n1058), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n728), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1079), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1056), .B1(new_n1083), .B2(G8), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT124), .B1(new_n1074), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(G8), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1056), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1050), .B1(new_n992), .B2(new_n1061), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(G288), .B2(new_n1069), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1073), .B1(new_n1090), .B2(new_n1067), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1039), .A2(KEYINPUT49), .A3(new_n1040), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(new_n1089), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT112), .B1(new_n1035), .B2(KEYINPUT49), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1041), .A2(new_n1037), .A3(new_n1042), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1093), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1091), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1088), .A2(new_n1097), .A3(new_n1098), .A4(new_n1065), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1085), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1966), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1081), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1028), .B1(new_n1001), .B2(KEYINPUT50), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1103), .A2(new_n768), .A3(new_n1063), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1050), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(new_n1104), .A3(G168), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(G8), .ZN(new_n1107));
  AOI21_X1  g682(.A(G168), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1108));
  OAI221_X1 g683(.A(KEYINPUT51), .B1(KEYINPUT121), .B2(new_n1105), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT51), .B1(new_n1105), .B2(KEYINPUT121), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1110), .A2(G8), .A3(new_n1106), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT62), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1080), .A2(new_n802), .A3(new_n992), .A4(new_n1058), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1057), .A2(KEYINPUT122), .A3(new_n802), .A4(new_n1058), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1117), .A3(KEYINPUT53), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1114), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(KEYINPUT123), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1103), .A2(new_n1063), .ZN(new_n1122));
  INV_X1    g697(.A(G1961), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT123), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1114), .A2(new_n1125), .A3(new_n1119), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1118), .A2(new_n1121), .A3(new_n1124), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(G171), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1109), .A2(new_n1130), .A3(new_n1111), .ZN(new_n1131));
  NAND4_X1  g706(.A1(new_n1100), .A2(new_n1113), .A3(new_n1129), .A4(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  AND2_X1   g708(.A1(new_n1105), .A2(G168), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n1088), .A2(new_n1097), .A3(new_n1065), .A4(new_n1134), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n1082), .B1(G2090), .B2(new_n1122), .ZN(new_n1136));
  OAI211_X1 g711(.A(KEYINPUT115), .B(new_n1049), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1136), .A2(G8), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1136), .B2(G8), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1105), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1139), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT113), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1091), .B2(new_n1096), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1045), .A2(KEYINPUT113), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  AOI22_X1  g721(.A1(new_n1133), .A2(new_n1135), .B1(new_n1142), .B2(new_n1146), .ZN(new_n1147));
  NOR3_X1   g722(.A1(new_n1096), .A2(G1976), .A3(G288), .ZN(new_n1148));
  NOR2_X1   g723(.A1(G305), .A2(G1981), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1089), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AND2_X1   g725(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(new_n1151), .B2(new_n1065), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1147), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1076), .A2(new_n1078), .A3(new_n1063), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(new_n759), .ZN(new_n1155));
  XNOR2_X1  g730(.A(KEYINPUT56), .B(G2072), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1080), .A2(new_n992), .A3(new_n1156), .A4(new_n1058), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT117), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND4_X1  g734(.A1(new_n1057), .A2(KEYINPUT117), .A3(new_n1156), .A4(new_n1058), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT116), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n1162), .A2(KEYINPUT57), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n571), .A2(new_n579), .A3(new_n580), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1162), .A2(KEYINPUT57), .ZN(new_n1165));
  XNOR2_X1  g740(.A(new_n1164), .B(new_n1165), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1155), .A2(new_n1161), .A3(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  AOI21_X1  g743(.A(new_n1166), .B1(new_n1155), .B2(new_n1161), .ZN(new_n1169));
  INV_X1    g744(.A(new_n1169), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1001), .A2(new_n1028), .A3(G2067), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1171), .B1(new_n1122), .B2(new_n667), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1172), .A2(new_n623), .ZN(new_n1173));
  AOI21_X1  g748(.A(new_n1168), .B1(new_n1170), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT119), .ZN(new_n1175));
  OAI21_X1  g750(.A(new_n1175), .B1(new_n621), .B2(new_n622), .ZN(new_n1176));
  INV_X1    g751(.A(KEYINPUT80), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n916), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n615), .A2(new_n620), .A3(KEYINPUT80), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1178), .A2(KEYINPUT119), .A3(new_n1179), .ZN(new_n1180));
  NAND4_X1  g755(.A1(new_n1176), .A2(new_n1180), .A3(KEYINPUT60), .A4(new_n1172), .ZN(new_n1181));
  OR2_X1    g756(.A1(new_n1172), .A2(KEYINPUT60), .ZN(new_n1182));
  INV_X1    g757(.A(new_n1171), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1060), .A2(new_n1063), .A3(new_n992), .ZN(new_n1184));
  OAI211_X1 g759(.A(KEYINPUT60), .B(new_n1183), .C1(new_n1184), .C2(G1348), .ZN(new_n1185));
  NAND3_X1  g760(.A1(new_n1185), .A2(KEYINPUT119), .A3(new_n623), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1181), .A2(new_n1182), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(KEYINPUT120), .ZN(new_n1188));
  INV_X1    g763(.A(KEYINPUT120), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1181), .A2(new_n1182), .A3(new_n1189), .A4(new_n1186), .ZN(new_n1190));
  AND2_X1   g765(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT118), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1001), .A2(new_n1028), .ZN(new_n1193));
  XNOR2_X1  g768(.A(KEYINPUT58), .B(G1341), .ZN(new_n1194));
  OAI22_X1  g769(.A1(new_n1081), .A2(G1996), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT59), .ZN(new_n1196));
  AND4_X1   g771(.A1(new_n1192), .A2(new_n1195), .A3(new_n562), .A4(new_n1196), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1192), .A2(new_n1196), .ZN(new_n1198));
  AOI22_X1  g773(.A1(new_n1195), .A2(new_n562), .B1(new_n1192), .B2(new_n1196), .ZN(new_n1199));
  NOR3_X1   g774(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(KEYINPUT61), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1201));
  INV_X1    g776(.A(KEYINPUT61), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n1170), .A2(new_n1202), .A3(new_n1167), .ZN(new_n1203));
  AOI21_X1  g778(.A(new_n1200), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(new_n1174), .B1(new_n1191), .B2(new_n1204), .ZN(new_n1205));
  AND2_X1   g780(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n1114), .A2(new_n1119), .ZN(new_n1207));
  NAND4_X1  g782(.A1(new_n1206), .A2(G301), .A3(new_n1121), .A4(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1128), .A2(new_n1208), .ZN(new_n1209));
  INV_X1    g784(.A(KEYINPUT54), .ZN(new_n1210));
  AOI22_X1  g785(.A1(new_n1209), .A2(new_n1210), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1211));
  OR2_X1    g786(.A1(new_n1127), .A2(G171), .ZN(new_n1212));
  AND3_X1   g787(.A1(new_n1206), .A2(new_n1121), .A3(new_n1207), .ZN(new_n1213));
  OAI211_X1 g788(.A(new_n1212), .B(KEYINPUT54), .C1(G301), .C2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1100), .A2(new_n1211), .A3(new_n1214), .ZN(new_n1215));
  OAI211_X1 g790(.A(new_n1132), .B(new_n1153), .C1(new_n1205), .C2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g791(.A1(G290), .A2(G1986), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1002), .B1(new_n1013), .B2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g793(.A1(new_n1022), .A2(new_n1218), .ZN(new_n1219));
  AND3_X1   g794(.A1(new_n1216), .A2(KEYINPUT125), .A3(new_n1219), .ZN(new_n1220));
  AOI21_X1  g795(.A(KEYINPUT125), .B1(new_n1216), .B2(new_n1219), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1027), .B1(new_n1220), .B2(new_n1221), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g797(.A(KEYINPUT127), .ZN(new_n1224));
  INV_X1    g798(.A(G319), .ZN(new_n1225));
  NOR2_X1   g799(.A1(G227), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g800(.A1(new_n712), .A2(new_n1226), .ZN(new_n1227));
  AOI21_X1  g801(.A(new_n1227), .B1(new_n678), .B2(new_n676), .ZN(new_n1228));
  AND2_X1   g802(.A1(new_n899), .A2(new_n1228), .ZN(new_n1229));
  AND3_X1   g803(.A1(new_n987), .A2(new_n1224), .A3(new_n1229), .ZN(new_n1230));
  AOI21_X1  g804(.A(new_n1224), .B1(new_n987), .B2(new_n1229), .ZN(new_n1231));
  NOR2_X1   g805(.A1(new_n1230), .A2(new_n1231), .ZN(G308));
  NAND2_X1  g806(.A1(new_n987), .A2(new_n1229), .ZN(new_n1233));
  NAND2_X1  g807(.A1(new_n1233), .A2(KEYINPUT127), .ZN(new_n1234));
  NAND3_X1  g808(.A1(new_n987), .A2(new_n1229), .A3(new_n1224), .ZN(new_n1235));
  NAND2_X1  g809(.A1(new_n1234), .A2(new_n1235), .ZN(G225));
endmodule


