//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1371,
    new_n1372, new_n1373;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NOR2_X1   g0011(.A1(G58), .A2(G68), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n206), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(KEYINPUT1), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  AND2_X1   g0024(.A1(new_n224), .A2(new_n208), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n211), .B(new_n218), .C1(new_n219), .C2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n225), .A2(new_n219), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT64), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n226), .A2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XOR2_X1   g0038(.A(G107), .B(G116), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g0040(.A(G50), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n241), .A2(G68), .ZN(new_n242));
  INV_X1    g0042(.A(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n240), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(G150), .ZN(new_n249));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  INV_X1    g0050(.A(new_n250), .ZN(new_n251));
  OAI22_X1  g0051(.A1(new_n249), .A2(new_n251), .B1(new_n201), .B2(new_n206), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n206), .A2(G33), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(KEYINPUT67), .ZN(new_n254));
  XOR2_X1   g0054(.A(KEYINPUT8), .B(G58), .Z(new_n255));
  AOI21_X1  g0055(.A(new_n252), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n216), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n262), .A2(new_n258), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n205), .A2(G20), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(G50), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n265), .B1(G50), .B2(new_n261), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT3), .B(G33), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G223), .ZN(new_n273));
  OAI22_X1  g0073(.A1(new_n272), .A2(new_n273), .B1(new_n202), .B2(new_n271), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT66), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n271), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G222), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n271), .A2(KEYINPUT66), .A3(G222), .A4(new_n276), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n274), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G33), .A2(G41), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G1), .A3(G13), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT65), .B(G41), .ZN(new_n285));
  INV_X1    g0085(.A(G45), .ZN(new_n286));
  AOI21_X1  g0086(.A(G1), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G274), .ZN(new_n288));
  INV_X1    g0088(.A(new_n216), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n288), .B1(new_n289), .B2(new_n282), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n205), .B1(G41), .B2(G45), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n283), .A2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n287), .A2(new_n290), .B1(new_n293), .B2(G226), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(G200), .B1(new_n284), .B2(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(G190), .B(new_n294), .C1(new_n281), .C2(new_n283), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n267), .A2(KEYINPUT9), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n270), .A2(new_n296), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n267), .B(new_n269), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n301), .A2(new_n302), .A3(new_n297), .A4(new_n296), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G169), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(new_n284), .B2(new_n295), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n307), .B(new_n294), .C1(new_n281), .C2(new_n283), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n268), .A3(new_n308), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n202), .B1(new_n205), .B2(G20), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n263), .A2(new_n310), .B1(new_n202), .B2(new_n262), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n255), .A2(new_n250), .B1(G20), .B2(G77), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT15), .B(G87), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n313), .B1(new_n253), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n312), .B1(new_n258), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n271), .A2(G232), .A3(new_n276), .ZN(new_n317));
  INV_X1    g0117(.A(G107), .ZN(new_n318));
  INV_X1    g0118(.A(G238), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n317), .B1(new_n318), .B2(new_n271), .C1(new_n272), .C2(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n283), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n287), .A2(new_n290), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n293), .A2(G244), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n322), .A2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n316), .B1(new_n327), .B2(new_n305), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n325), .B1(new_n321), .B2(new_n320), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(new_n307), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n327), .A2(G200), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n315), .A2(new_n258), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n311), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n334), .B1(new_n329), .B2(G190), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n331), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n304), .A2(new_n309), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT68), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT68), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n304), .A2(new_n336), .A3(new_n339), .A4(new_n309), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT77), .ZN(new_n342));
  INV_X1    g0142(.A(G33), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT3), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT3), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(G33), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n344), .A2(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT7), .B1(new_n347), .B2(new_n206), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT7), .ZN(new_n349));
  AOI211_X1 g0149(.A(new_n349), .B(G20), .C1(new_n344), .C2(new_n346), .ZN(new_n350));
  OAI21_X1  g0150(.A(G68), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  AND2_X1   g0151(.A1(G58), .A2(G68), .ZN(new_n352));
  OAI21_X1  g0152(.A(G20), .B1(new_n352), .B2(new_n212), .ZN(new_n353));
  INV_X1    g0153(.A(G159), .ZN(new_n354));
  NOR4_X1   g0154(.A1(new_n354), .A2(KEYINPUT72), .A3(G20), .A4(G33), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT72), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n356), .B1(new_n250), .B2(G159), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n353), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT73), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT73), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n360), .B(new_n353), .C1(new_n355), .C2(new_n357), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n351), .A2(KEYINPUT16), .A3(new_n359), .A4(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT74), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n349), .B1(new_n271), .B2(G20), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n347), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n206), .A2(new_n343), .A3(G159), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT72), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n250), .A2(new_n356), .A3(G159), .ZN(new_n370));
  XNOR2_X1  g0170(.A(G58), .B(G68), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n369), .A2(new_n370), .B1(new_n371), .B2(G20), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n367), .A2(G68), .B1(new_n372), .B2(new_n360), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n373), .A2(KEYINPUT74), .A3(KEYINPUT16), .A4(new_n359), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n364), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT16), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n243), .B1(new_n365), .B2(new_n366), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n376), .B1(new_n377), .B2(new_n358), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n258), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n375), .A2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(G200), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n271), .A2(G226), .A3(G1698), .ZN(new_n383));
  NAND2_X1  g0183(.A1(G33), .A2(G87), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n383), .B(new_n384), .C1(new_n277), .C2(new_n273), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n385), .A2(new_n321), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n287), .A2(new_n290), .B1(new_n293), .B2(G232), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n382), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n386), .A2(new_n387), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n388), .B1(new_n390), .B2(G190), .ZN(new_n391));
  INV_X1    g0191(.A(new_n263), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n255), .A2(new_n264), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n392), .A2(new_n393), .B1(new_n261), .B2(new_n255), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n394), .B(KEYINPUT75), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n381), .A2(new_n391), .A3(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT17), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n379), .B1(new_n364), .B2(new_n374), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(new_n395), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(KEYINPUT17), .A3(new_n391), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n389), .A2(G169), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n403), .B1(new_n307), .B2(new_n389), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n400), .B2(new_n395), .ZN(new_n405));
  NOR2_X1   g0205(.A1(KEYINPUT76), .A2(KEYINPUT18), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n399), .A2(new_n402), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT76), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n405), .A2(KEYINPUT18), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT18), .ZN(new_n411));
  OAI211_X1 g0211(.A(new_n404), .B(new_n411), .C1(new_n400), .C2(new_n395), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n409), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n271), .A2(G232), .A3(G1698), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G97), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n344), .A2(new_n346), .A3(G226), .A4(new_n276), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT69), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n271), .A2(KEYINPUT69), .A3(G226), .A4(new_n276), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n283), .B1(new_n417), .B2(new_n422), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n287), .A2(new_n290), .B1(new_n293), .B2(G238), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT13), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT13), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n415), .A2(new_n416), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n428), .B1(new_n420), .B2(new_n421), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n427), .B(new_n424), .C1(new_n429), .C2(new_n283), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(G169), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT14), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n433), .A2(KEYINPUT71), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT70), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n426), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g0237(.A(KEYINPUT70), .B(KEYINPUT13), .C1(new_n423), .C2(new_n425), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n437), .A2(G179), .A3(new_n438), .A4(new_n430), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n431), .B(G169), .C1(KEYINPUT71), .C2(new_n433), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n254), .A2(G77), .ZN(new_n442));
  AOI22_X1  g0242(.A1(new_n250), .A2(G50), .B1(G20), .B2(new_n243), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n259), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  OR2_X1    g0244(.A1(new_n444), .A2(KEYINPUT11), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n444), .A2(KEYINPUT11), .ZN(new_n446));
  OAI21_X1  g0246(.A(KEYINPUT12), .B1(new_n261), .B2(G68), .ZN(new_n447));
  OR3_X1    g0247(.A1(new_n261), .A2(KEYINPUT12), .A3(G68), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n243), .B1(new_n205), .B2(G20), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n447), .A2(new_n448), .B1(new_n263), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n445), .A2(new_n446), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n441), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n451), .B1(new_n431), .B2(G200), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n437), .A2(G190), .A3(new_n438), .A4(new_n430), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n341), .A2(new_n342), .A3(new_n414), .A4(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n457), .A2(new_n338), .A3(new_n340), .ZN(new_n459));
  INV_X1    g0259(.A(new_n414), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT77), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n463));
  AND2_X1   g0263(.A1(new_n463), .A2(new_n206), .ZN(new_n464));
  INV_X1    g0264(.A(G87), .ZN(new_n465));
  INV_X1    g0265(.A(G97), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n465), .A2(new_n466), .A3(new_n318), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT79), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n465), .A2(new_n466), .A3(new_n318), .A4(KEYINPUT79), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n344), .A2(new_n346), .A3(new_n206), .A4(G68), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT19), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n473), .B1(new_n253), .B2(new_n466), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n258), .B1(new_n471), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n314), .A2(new_n262), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n343), .A2(G1), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n262), .A2(new_n258), .A3(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n314), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n476), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(G250), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n483), .B1(new_n286), .B2(G1), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n205), .A2(new_n288), .A3(G45), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n283), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n344), .A2(new_n346), .A3(G244), .A4(G1698), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n344), .A2(new_n346), .A3(G238), .A4(new_n276), .ZN(new_n489));
  NAND2_X1  g0289(.A1(G33), .A2(G116), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n487), .B1(new_n491), .B2(new_n321), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n307), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n482), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n491), .A2(new_n321), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n486), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n305), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n479), .A2(G87), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n476), .A2(new_n477), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(G190), .ZN(new_n500));
  AOI211_X1 g0300(.A(new_n500), .B(new_n487), .C1(new_n491), .C2(new_n321), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n496), .A2(G200), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n494), .A2(new_n497), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n344), .A2(new_n346), .A3(new_n206), .A4(G87), .ZN(new_n505));
  NAND2_X1  g0305(.A1(KEYINPUT80), .A2(KEYINPUT22), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n505), .A2(new_n507), .ZN(new_n508));
  NAND4_X1  g0308(.A1(new_n271), .A2(new_n206), .A3(G87), .A4(new_n506), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(KEYINPUT82), .A2(KEYINPUT24), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT81), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(new_n490), .B2(G20), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n206), .A2(KEYINPUT81), .A3(G33), .A4(G116), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  OAI21_X1  g0315(.A(KEYINPUT23), .B1(new_n206), .B2(G107), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT23), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n517), .A2(new_n318), .A3(G20), .ZN(new_n518));
  NAND2_X1  g0318(.A1(KEYINPUT82), .A2(KEYINPUT24), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n516), .A2(new_n518), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n515), .A2(new_n520), .ZN(new_n521));
  AND3_X1   g0321(.A1(new_n510), .A2(new_n511), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n511), .B1(new_n510), .B2(new_n521), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n258), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT83), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT25), .ZN(new_n526));
  AOI211_X1 g0326(.A(G107), .B(new_n261), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n525), .A2(new_n526), .ZN(new_n528));
  OR2_X1    g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n528), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n529), .A2(new_n530), .B1(G107), .B2(new_n479), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n524), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(G41), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(KEYINPUT65), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT65), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G41), .ZN(new_n536));
  AOI21_X1  g0336(.A(KEYINPUT5), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT5), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n205), .B(G45), .C1(new_n538), .C2(G41), .ZN(new_n539));
  OAI211_X1 g0339(.A(G264), .B(new_n283), .C1(new_n537), .C2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n538), .A2(G41), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n205), .A2(G45), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n290), .B(new_n543), .C1(KEYINPUT5), .C2(new_n285), .ZN(new_n544));
  INV_X1    g0344(.A(G294), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n343), .A2(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(G250), .A2(G1698), .ZN(new_n547));
  INV_X1    g0347(.A(G257), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n547), .B1(new_n548), .B2(G1698), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n546), .B1(new_n549), .B2(new_n271), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n540), .B(new_n544), .C1(new_n283), .C2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(new_n305), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(G1698), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(G250), .B2(G1698), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n554), .A2(new_n347), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n321), .B1(new_n555), .B2(new_n546), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n556), .A2(new_n307), .A3(new_n544), .A4(new_n540), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n552), .A2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n532), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n551), .A2(new_n382), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n556), .A2(new_n500), .A3(new_n544), .A4(new_n540), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(new_n524), .A3(new_n531), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n504), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  NAND4_X1  g0365(.A1(new_n344), .A2(new_n346), .A3(G244), .A4(new_n276), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT4), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G33), .A2(G283), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(G250), .A2(G1698), .ZN(new_n571));
  NAND2_X1  g0371(.A1(KEYINPUT4), .A2(G244), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n571), .B1(new_n572), .B2(G1698), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n570), .B1(new_n271), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(KEYINPUT78), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT78), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n568), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n321), .A3(new_n578), .ZN(new_n579));
  OAI211_X1 g0379(.A(G257), .B(new_n283), .C1(new_n537), .C2(new_n539), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n544), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n307), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT6), .ZN(new_n584));
  NOR3_X1   g0384(.A1(new_n584), .A2(new_n466), .A3(G107), .ZN(new_n585));
  XNOR2_X1  g0385(.A(G97), .B(G107), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n585), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  OAI22_X1  g0387(.A1(new_n587), .A2(new_n206), .B1(new_n202), .B2(new_n251), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n318), .B1(new_n365), .B2(new_n366), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n258), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n262), .A2(new_n466), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n479), .A2(G97), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n283), .B1(new_n575), .B2(KEYINPUT78), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n581), .B1(new_n594), .B2(new_n578), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n583), .B(new_n593), .C1(G169), .C2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n579), .A2(G190), .A3(new_n582), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n592), .A2(new_n591), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n367), .A2(G107), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n251), .A2(new_n202), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n586), .A2(new_n584), .ZN(new_n601));
  INV_X1    g0401(.A(new_n585), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n600), .B1(new_n603), .B2(G20), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n598), .B1(new_n605), .B2(new_n258), .ZN(new_n606));
  OAI211_X1 g0406(.A(new_n597), .B(new_n606), .C1(new_n382), .C2(new_n595), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n596), .A2(new_n607), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n569), .B(new_n206), .C1(G33), .C2(new_n466), .ZN(new_n609));
  INV_X1    g0409(.A(G116), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(G20), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n609), .A2(new_n258), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT20), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n609), .A2(KEYINPUT20), .A3(new_n258), .A4(new_n611), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n261), .A2(G116), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(new_n479), .B2(G116), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(G270), .B(new_n283), .C1(new_n537), .C2(new_n539), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n621), .A2(new_n544), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n344), .A2(new_n346), .A3(G264), .A4(G1698), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n344), .A2(new_n346), .A3(G257), .A4(new_n276), .ZN(new_n624));
  INV_X1    g0424(.A(G303), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n271), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n321), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n622), .A2(G190), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n544), .A3(new_n621), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n620), .B(new_n628), .C1(new_n630), .C2(new_n382), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(G179), .A3(new_n619), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n305), .B1(new_n616), .B2(new_n618), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT21), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n633), .A2(new_n634), .A3(new_n629), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n634), .B1(new_n633), .B2(new_n629), .ZN(new_n636));
  OAI211_X1 g0436(.A(new_n631), .B(new_n632), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n565), .A2(new_n608), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n462), .A2(new_n638), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n639), .B(KEYINPUT84), .ZN(G372));
  INV_X1    g0440(.A(new_n309), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n454), .A2(new_n455), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n453), .B1(new_n642), .B2(new_n331), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n399), .A2(new_n402), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n410), .B(new_n412), .C1(new_n643), .C2(new_n644), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n641), .B1(new_n645), .B2(new_n304), .ZN(new_n646));
  INV_X1    g0446(.A(new_n462), .ZN(new_n647));
  AND3_X1   g0447(.A1(new_n476), .A2(new_n477), .A3(new_n498), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n491), .A2(new_n321), .ZN(new_n649));
  XNOR2_X1  g0449(.A(new_n486), .B(KEYINPUT85), .ZN(new_n650));
  OAI21_X1  g0450(.A(G200), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT86), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n648), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT85), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n486), .B(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n382), .B1(new_n655), .B2(new_n495), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT86), .B1(new_n656), .B2(new_n499), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n492), .A2(G190), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n653), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n655), .A2(new_n495), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(new_n305), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n494), .A2(new_n661), .ZN(new_n662));
  AND3_X1   g0462(.A1(new_n659), .A2(new_n564), .A3(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT87), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n596), .A2(new_n607), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n620), .A2(new_n629), .A3(new_n307), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n633), .A2(new_n629), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(KEYINPUT21), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n633), .A2(new_n634), .A3(new_n629), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n560), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n659), .A2(new_n564), .A3(new_n662), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT87), .B1(new_n673), .B2(new_n608), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n666), .A2(new_n672), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n596), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n676), .A2(new_n677), .A3(new_n662), .A4(new_n659), .ZN(new_n678));
  XNOR2_X1  g0478(.A(new_n662), .B(KEYINPUT88), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n648), .A2(new_n503), .A3(new_n658), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n497), .A2(new_n482), .A3(new_n493), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(KEYINPUT26), .B1(new_n596), .B2(new_n682), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n678), .A2(new_n679), .A3(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n675), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n646), .B1(new_n647), .B2(new_n686), .ZN(G369));
  NAND3_X1  g0487(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(G343), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n671), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT90), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n532), .A2(new_n694), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n560), .A2(new_n697), .A3(new_n564), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n560), .B2(new_n693), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n558), .B1(new_n524), .B2(new_n531), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n700), .B1(new_n701), .B2(new_n693), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n694), .A2(new_n619), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(KEYINPUT89), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n706), .B1(new_n637), .B2(new_n705), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n703), .A2(KEYINPUT89), .A3(new_n705), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(G330), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(new_n699), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n702), .A2(new_n712), .ZN(G399));
  INV_X1    g0513(.A(new_n209), .ZN(new_n714));
  INV_X1    g0514(.A(new_n285), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n205), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n469), .A2(new_n470), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n610), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI22_X1  g0520(.A1(new_n717), .A2(new_n720), .B1(new_n215), .B2(new_n716), .ZN(new_n721));
  XOR2_X1   g0521(.A(new_n721), .B(KEYINPUT28), .Z(new_n722));
  NOR3_X1   g0522(.A1(new_n686), .A2(KEYINPUT29), .A3(new_n694), .ZN(new_n723));
  INV_X1    g0523(.A(KEYINPUT29), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n608), .A2(KEYINPUT94), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT94), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n596), .A2(new_n607), .A3(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n725), .A2(new_n663), .A3(new_n672), .A4(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(KEYINPUT95), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n703), .A2(new_n701), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(new_n673), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT95), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n731), .A2(new_n732), .A3(new_n725), .A4(new_n727), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n659), .A2(new_n662), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n734), .A2(KEYINPUT26), .A3(new_n676), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n677), .B1(new_n596), .B2(new_n682), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT93), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  OAI211_X1 g0538(.A(KEYINPUT93), .B(new_n677), .C1(new_n596), .C2(new_n682), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n735), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n729), .A2(new_n679), .A3(new_n733), .A4(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n724), .B1(new_n741), .B2(new_n693), .ZN(new_n742));
  INV_X1    g0542(.A(new_n564), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n743), .A2(new_n701), .A3(new_n682), .ZN(new_n744));
  INV_X1    g0544(.A(new_n637), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n744), .A2(new_n665), .A3(new_n745), .A4(new_n693), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(KEYINPUT31), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n556), .A2(G179), .A3(new_n540), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n749), .A2(new_n492), .A3(new_n627), .A4(new_n622), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n579), .A2(new_n582), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n748), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AND2_X1   g0552(.A1(new_n551), .A2(new_n307), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n751), .A2(new_n753), .A3(new_n629), .A4(new_n660), .ZN(new_n754));
  AND4_X1   g0554(.A1(G179), .A2(new_n492), .A3(new_n540), .A4(new_n556), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n755), .A2(new_n595), .A3(KEYINPUT30), .A4(new_n630), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n752), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT92), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n752), .A2(new_n756), .A3(KEYINPUT92), .A4(new_n754), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n759), .A2(new_n694), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n747), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n752), .A2(new_n754), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(KEYINPUT91), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(new_n756), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n763), .A2(KEYINPUT91), .ZN(new_n766));
  OAI211_X1 g0566(.A(KEYINPUT31), .B(new_n694), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n710), .B1(new_n762), .B2(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n723), .A2(new_n742), .A3(new_n768), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n722), .B1(new_n769), .B2(G1), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT96), .ZN(G364));
  NAND2_X1  g0571(.A1(new_n206), .A2(G13), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT97), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(G45), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n717), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n711), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n709), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n777), .B1(G330), .B2(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G13), .A2(G33), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n781), .A2(G20), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n209), .A2(G355), .A3(new_n271), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n714), .A2(new_n271), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(G45), .B2(new_n214), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n247), .A2(new_n286), .ZN(new_n788));
  OAI221_X1 g0588(.A(new_n785), .B1(G116), .B2(new_n209), .C1(new_n787), .C2(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n216), .B1(G20), .B2(new_n305), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n782), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n775), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g0592(.A(KEYINPUT99), .B1(new_n307), .B2(G200), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n206), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n307), .A2(KEYINPUT99), .A3(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(G190), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n797), .A2(G283), .ZN(new_n798));
  NAND2_X1  g0598(.A1(G20), .A2(G179), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT98), .Z(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G200), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n500), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G326), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n796), .A2(new_n500), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n803), .B1(new_n625), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n801), .A2(G190), .ZN(new_n807));
  XNOR2_X1  g0607(.A(KEYINPUT33), .B(G317), .ZN(new_n808));
  AOI211_X1 g0608(.A(new_n798), .B(new_n806), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G190), .A2(G200), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n810), .A2(G20), .A3(new_n307), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n271), .B1(new_n812), .B2(G329), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n500), .A2(G179), .A3(G200), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n206), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n500), .A2(G200), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n800), .A2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G322), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n813), .B1(new_n545), .B2(new_n815), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n800), .A2(new_n810), .ZN(new_n820));
  INV_X1    g0620(.A(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n819), .B1(G311), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n815), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(G97), .ZN(new_n824));
  INV_X1    g0624(.A(new_n807), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n825), .B2(new_n243), .ZN(new_n826));
  XNOR2_X1  g0626(.A(new_n826), .B(KEYINPUT100), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n804), .A2(G87), .ZN(new_n828));
  INV_X1    g0628(.A(new_n797), .ZN(new_n829));
  INV_X1    g0629(.A(new_n802), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n828), .B1(new_n829), .B2(new_n318), .C1(new_n830), .C2(new_n241), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n812), .A2(G159), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n347), .B1(new_n832), .B2(KEYINPUT32), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(KEYINPUT32), .B2(new_n832), .ZN(new_n834));
  INV_X1    g0634(.A(G58), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n835), .A2(new_n817), .B1(new_n820), .B2(new_n202), .ZN(new_n836));
  NOR3_X1   g0636(.A1(new_n831), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n809), .A2(new_n822), .B1(new_n827), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n790), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n792), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n779), .B1(new_n784), .B2(new_n840), .ZN(G396));
  NAND2_X1  g0641(.A1(new_n329), .A2(G190), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n332), .A2(new_n842), .A3(new_n316), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n334), .A2(new_n694), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n843), .A2(new_n844), .B1(new_n328), .B2(new_n330), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n328), .A2(new_n330), .A3(new_n693), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  OAI21_X1  g0647(.A(KEYINPUT102), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT102), .ZN(new_n849));
  AOI22_X1  g0649(.A1(new_n335), .A2(new_n332), .B1(new_n334), .B2(new_n694), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n849), .B(new_n846), .C1(new_n850), .C2(new_n331), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n686), .B2(new_n694), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n848), .A2(new_n851), .A3(new_n693), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n685), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n768), .B1(new_n853), .B2(new_n856), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(new_n717), .B2(new_n774), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n853), .A2(new_n768), .A3(new_n856), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n790), .A2(new_n780), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n775), .B1(new_n202), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n271), .B1(new_n812), .B2(G311), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n824), .B(new_n863), .C1(new_n817), .C2(new_n545), .ZN(new_n864));
  XOR2_X1   g0664(.A(KEYINPUT101), .B(G283), .Z(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  AOI22_X1  g0666(.A1(G303), .A2(new_n802), .B1(new_n807), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n797), .A2(G87), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n867), .B(new_n868), .C1(new_n318), .C2(new_n805), .ZN(new_n869));
  AOI211_X1 g0669(.A(new_n864), .B(new_n869), .C1(G116), .C2(new_n821), .ZN(new_n870));
  INV_X1    g0670(.A(new_n817), .ZN(new_n871));
  AOI22_X1  g0671(.A1(G143), .A2(new_n871), .B1(new_n821), .B2(G159), .ZN(new_n872));
  INV_X1    g0672(.A(G137), .ZN(new_n873));
  OAI221_X1 g0673(.A(new_n872), .B1(new_n825), .B2(new_n249), .C1(new_n873), .C2(new_n830), .ZN(new_n874));
  XNOR2_X1  g0674(.A(new_n874), .B(KEYINPUT34), .ZN(new_n875));
  INV_X1    g0675(.A(G132), .ZN(new_n876));
  OAI221_X1 g0676(.A(new_n271), .B1(new_n876), .B2(new_n811), .C1(new_n815), .C2(new_n835), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n829), .A2(new_n243), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n877), .B(new_n878), .C1(G50), .C2(new_n804), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n870), .B1(new_n875), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n852), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n862), .B1(new_n880), .B2(new_n839), .C1(new_n881), .C2(new_n781), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n860), .A2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(G384));
  OR2_X1    g0684(.A1(new_n603), .A2(KEYINPUT35), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n603), .A2(KEYINPUT35), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n885), .A2(G116), .A3(new_n217), .A4(new_n886), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT36), .Z(new_n888));
  OR3_X1    g0688(.A1(new_n214), .A2(new_n202), .A3(new_n352), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n205), .B(G13), .C1(new_n889), .C2(new_n242), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n693), .B1(new_n757), .B2(new_n758), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n746), .A2(KEYINPUT31), .B1(new_n760), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n892), .A2(KEYINPUT31), .A3(new_n760), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(KEYINPUT104), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT104), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT31), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(new_n638), .B2(new_n693), .ZN(new_n899));
  INV_X1    g0699(.A(new_n761), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n897), .B(new_n894), .C1(new_n899), .C2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n896), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n462), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n903), .B(KEYINPUT105), .Z(new_n904));
  OAI21_X1  g0704(.A(new_n692), .B1(new_n400), .B2(new_n395), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n410), .A2(new_n412), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n906), .B1(new_n644), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n397), .A2(new_n405), .A3(new_n905), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT37), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT37), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n397), .A2(new_n405), .A3(new_n905), .A4(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n908), .A2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT38), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n373), .A2(new_n359), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n259), .B1(new_n917), .B2(new_n376), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n375), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(new_n394), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n691), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n408), .B2(new_n413), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n389), .A2(G200), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n500), .B2(new_n389), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n400), .A2(new_n924), .A3(new_n395), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n390), .A2(G179), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n919), .A2(new_n920), .B1(new_n403), .B2(new_n926), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n925), .A2(new_n927), .A3(new_n921), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n912), .B1(new_n928), .B2(new_n911), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n922), .A2(new_n929), .A3(KEYINPUT38), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n916), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n451), .A2(new_n694), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n452), .A2(new_n642), .A3(new_n932), .ZN(new_n933));
  OAI211_X1 g0733(.A(new_n451), .B(new_n694), .C1(new_n456), .C2(new_n441), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n881), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n931), .A2(new_n902), .A3(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT40), .ZN(new_n939));
  INV_X1    g0739(.A(new_n921), .ZN(new_n940));
  AND3_X1   g0740(.A1(new_n399), .A2(new_n402), .A3(new_n407), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n907), .A2(KEYINPUT76), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n912), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n919), .A2(new_n920), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n404), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n940), .A2(new_n946), .A3(new_n397), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n944), .B1(KEYINPUT37), .B2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n915), .B1(new_n943), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(KEYINPUT40), .B1(new_n949), .B2(new_n930), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n936), .B1(new_n901), .B2(new_n896), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n939), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n904), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n904), .A2(new_n953), .ZN(new_n955));
  NOR3_X1   g0755(.A1(new_n954), .A2(new_n955), .A3(new_n710), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT103), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n856), .A2(new_n957), .A3(new_n846), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n854), .B1(new_n675), .B2(new_n684), .ZN(new_n959));
  OAI21_X1  g0759(.A(KEYINPUT103), .B1(new_n959), .B2(new_n847), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n949), .A2(new_n930), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n961), .A2(new_n962), .A3(new_n935), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT39), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n931), .A2(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n452), .A2(new_n694), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n949), .A2(KEYINPUT39), .A3(new_n930), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n907), .A2(new_n691), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n963), .A2(new_n968), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n462), .B1(new_n742), .B2(new_n723), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n646), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n970), .B(new_n972), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n956), .A2(new_n973), .B1(new_n205), .B2(new_n773), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n956), .A2(new_n973), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n891), .B1(new_n974), .B2(new_n975), .ZN(G367));
  INV_X1    g0776(.A(new_n786), .ZN(new_n977));
  OAI221_X1 g0777(.A(new_n791), .B1(new_n209), .B2(new_n314), .C1(new_n977), .C2(new_n236), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n776), .ZN(new_n979));
  XOR2_X1   g0779(.A(new_n979), .B(KEYINPUT109), .Z(new_n980));
  NAND2_X1  g0780(.A1(new_n694), .A2(new_n499), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n679), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n734), .A2(new_n981), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n802), .A2(G311), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n807), .A2(G294), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n797), .A2(G97), .ZN(new_n987));
  AND3_X1   g0787(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n271), .B1(new_n812), .B2(G317), .ZN(new_n989));
  OAI221_X1 g0789(.A(new_n989), .B1(new_n318), .B2(new_n815), .C1(new_n817), .C2(new_n625), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(new_n821), .B2(new_n866), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n804), .A2(G116), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT46), .ZN(new_n993));
  NAND3_X1  g0793(.A1(new_n988), .A2(new_n991), .A3(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT110), .Z(new_n995));
  NAND2_X1  g0795(.A1(new_n797), .A2(G77), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n805), .B2(new_n835), .C1(new_n825), .C2(new_n354), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n823), .A2(G68), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n817), .B2(new_n249), .ZN(new_n999));
  INV_X1    g0799(.A(KEYINPUT111), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n802), .A2(G143), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n271), .B1(new_n811), .B2(new_n873), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(new_n821), .B2(G50), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n999), .A2(new_n1000), .ZN(new_n1006));
  NOR3_X1   g0806(.A1(new_n997), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n995), .A2(new_n1007), .ZN(new_n1008));
  AND2_X1   g0808(.A1(new_n1008), .A2(KEYINPUT47), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n790), .B1(new_n1008), .B2(KEYINPUT47), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n980), .B1(new_n783), .B2(new_n984), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  OAI211_X1 g0811(.A(new_n725), .B(new_n727), .C1(new_n606), .C2(new_n693), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n596), .B2(new_n693), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n700), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n596), .B1(new_n1012), .B2(new_n560), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1014), .A2(KEYINPUT42), .B1(new_n693), .B2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(KEYINPUT42), .B2(new_n1014), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT43), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n984), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1017), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT106), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1019), .A2(new_n1018), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n711), .A2(new_n699), .A3(new_n1013), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1023), .B(new_n1024), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n774), .A2(G1), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n702), .A2(new_n1013), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT45), .Z(new_n1028));
  NOR2_X1   g0828(.A1(new_n702), .A2(new_n1013), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT44), .ZN(new_n1030));
  AND3_X1   g0830(.A1(new_n1028), .A2(new_n712), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n712), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1032));
  NOR2_X1   g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n696), .B(new_n699), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n711), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1034), .B1(KEYINPUT107), .B2(new_n1035), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n711), .B(KEYINPUT107), .Z(new_n1037));
  AOI21_X1  g0837(.A(new_n1036), .B1(new_n1037), .B2(new_n1034), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1038), .A2(KEYINPUT108), .A3(new_n769), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n769), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT108), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1033), .A2(new_n1039), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n769), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n716), .B(KEYINPUT41), .Z(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1026), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1011), .B1(new_n1025), .B2(new_n1047), .ZN(G387));
  OR2_X1    g0848(.A1(new_n699), .A2(new_n783), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n786), .B1(new_n233), .B2(new_n286), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n719), .A2(new_n209), .A3(new_n271), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n255), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n1054));
  OR3_X1    g0854(.A1(new_n1053), .A2(new_n1054), .A3(G50), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1054), .B1(new_n1053), .B2(G50), .ZN(new_n1056));
  AOI21_X1  g0856(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n720), .A2(new_n1055), .A3(new_n1056), .A4(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1052), .A2(new_n1058), .B1(new_n318), .B2(new_n714), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n791), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n776), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n823), .A2(new_n480), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n347), .B1(new_n812), .B2(G150), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(new_n817), .C2(new_n241), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1064), .B1(G68), .B2(new_n821), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G159), .A2(new_n802), .B1(new_n807), .B2(new_n255), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n804), .A2(G77), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1065), .A2(new_n1066), .A3(new_n987), .A4(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n271), .B1(new_n812), .B2(G326), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n805), .A2(new_n545), .B1(new_n815), .B2(new_n865), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G303), .A2(new_n821), .B1(new_n871), .B2(G317), .ZN(new_n1071));
  INV_X1    g0871(.A(G311), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1071), .B1(new_n825), .B2(new_n1072), .C1(new_n818), .C2(new_n830), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT48), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1070), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1075), .B1(new_n1074), .B2(new_n1073), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT49), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1069), .B1(new_n610), .B2(new_n829), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1068), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1061), .B1(new_n1080), .B2(new_n790), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n1038), .A2(new_n1026), .B1(new_n1049), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1040), .A2(new_n716), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1038), .A2(new_n769), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(G393));
  INV_X1    g0885(.A(new_n716), .ZN(new_n1086));
  OR2_X1    g0886(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1086), .B1(new_n1087), .B2(new_n1040), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n1043), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n786), .A2(new_n240), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1060), .B1(G97), .B2(new_n714), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n775), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n271), .B1(new_n812), .B2(G322), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n610), .B2(new_n815), .C1(new_n820), .C2(new_n545), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n825), .A2(new_n625), .B1(new_n805), .B2(new_n865), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n1094), .B(new_n1095), .C1(G107), .C2(new_n797), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n802), .A2(G317), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n1072), .B2(new_n817), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT52), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n830), .A2(new_n249), .B1(new_n817), .B2(new_n354), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT51), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n807), .A2(G50), .B1(new_n821), .B2(new_n255), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1102), .A2(KEYINPUT113), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1102), .A2(KEYINPUT113), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n804), .A2(G68), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n823), .A2(G77), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n347), .B1(new_n812), .B2(G143), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n868), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  NOR3_X1   g0908(.A1(new_n1103), .A2(new_n1104), .A3(new_n1108), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1096), .A2(new_n1099), .B1(new_n1101), .B2(new_n1109), .ZN(new_n1110));
  OAI221_X1 g0910(.A(new_n1092), .B1(new_n839), .B2(new_n1110), .C1(new_n1013), .C2(new_n783), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1026), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1111), .B1(new_n1087), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1089), .A2(new_n1114), .ZN(G390));
  NAND3_X1  g0915(.A1(new_n768), .A2(new_n881), .A3(new_n935), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n933), .A2(new_n934), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(new_n958), .B2(new_n960), .ZN(new_n1118));
  AND3_X1   g0918(.A1(new_n949), .A2(KEYINPUT39), .A3(new_n930), .ZN(new_n1119));
  AOI21_X1  g0919(.A(KEYINPUT39), .B1(new_n916), .B2(new_n930), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n1118), .A2(new_n966), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n741), .A2(new_n693), .A3(new_n881), .ZN(new_n1122));
  AND3_X1   g0922(.A1(new_n1122), .A2(KEYINPUT114), .A3(new_n846), .ZN(new_n1123));
  AOI21_X1  g0923(.A(KEYINPUT114), .B1(new_n1122), .B2(new_n846), .ZN(new_n1124));
  NOR3_X1   g0924(.A1(new_n1123), .A2(new_n1124), .A3(new_n1117), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n966), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n931), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1116), .B(new_n1121), .C1(new_n1125), .C2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1122), .A2(new_n846), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT114), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1122), .A2(KEYINPUT114), .A3(new_n846), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1131), .A2(new_n935), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1127), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n957), .B1(new_n856), .B2(new_n846), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n959), .A2(KEYINPUT103), .A3(new_n847), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n935), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n1126), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n965), .A2(new_n967), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n1133), .A2(new_n1134), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n902), .A2(G330), .A3(new_n937), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1128), .B(new_n1026), .C1(new_n1140), .C2(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT118), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1139), .A2(new_n780), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n775), .B1(new_n1053), .B2(new_n861), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n271), .B1(new_n812), .B2(G294), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1106), .B(new_n1146), .C1(new_n817), .C2(new_n610), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(G107), .A2(new_n807), .B1(new_n802), .B2(G283), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n878), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n1149), .A3(new_n828), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1147), .B(new_n1150), .C1(G97), .C2(new_n821), .ZN(new_n1151));
  OR2_X1    g0951(.A1(new_n1151), .A2(KEYINPUT117), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(KEYINPUT117), .ZN(new_n1153));
  OAI22_X1  g0953(.A1(new_n825), .A2(new_n873), .B1(new_n829), .B2(new_n241), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1154), .B1(G128), .B2(new_n802), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n804), .A2(G150), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT53), .Z(new_n1157));
  AOI21_X1  g0957(.A(new_n347), .B1(new_n812), .B2(G125), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(KEYINPUT54), .B(G143), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1158), .B1(new_n354), .B2(new_n815), .C1(new_n820), .C2(new_n1159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G132), .B2(new_n871), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1155), .A2(new_n1157), .A3(new_n1161), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1152), .A2(new_n1153), .A3(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n1144), .B(new_n1145), .C1(new_n839), .C2(new_n1163), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n1142), .A2(new_n1143), .A3(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1143), .B1(new_n1142), .B2(new_n1164), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT116), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n902), .A2(G330), .A3(new_n881), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1169), .A2(new_n1117), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(KEYINPUT115), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1116), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT115), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1169), .A2(new_n1174), .A3(new_n1117), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1171), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n768), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1117), .B1(new_n1177), .B2(new_n852), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n1141), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n961), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n462), .A2(G330), .A3(new_n902), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n971), .A2(new_n1182), .A3(new_n646), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1128), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1168), .B(new_n716), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1183), .B1(new_n1176), .B2(new_n1180), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1190), .B(new_n1128), .C1(new_n1141), .C2(new_n1140), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1168), .B1(new_n1191), .B2(new_n716), .ZN(new_n1192));
  OAI21_X1  g0992(.A(new_n1167), .B1(new_n1189), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(KEYINPUT119), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT119), .ZN(new_n1195));
  OAI211_X1 g0995(.A(new_n1167), .B(new_n1195), .C1(new_n1189), .C2(new_n1192), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1194), .A2(new_n1196), .ZN(G378));
  NAND2_X1  g0997(.A1(new_n304), .A2(new_n309), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n268), .A2(new_n692), .ZN(new_n1199));
  XNOR2_X1  g0999(.A(new_n1198), .B(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1200), .B(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1203), .A2(new_n780), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n241), .B1(G33), .B2(G41), .C1(new_n715), .C2(new_n271), .ZN(new_n1205));
  AOI211_X1 g1005(.A(new_n271), .B(new_n715), .C1(G283), .C2(new_n812), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1206), .A2(new_n998), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n318), .B2(new_n817), .C1(new_n314), .C2(new_n820), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1067), .B1(new_n829), .B2(new_n835), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n466), .A2(new_n825), .B1(new_n830), .B2(new_n610), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  XOR2_X1   g1011(.A(KEYINPUT120), .B(KEYINPUT58), .Z(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1205), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT121), .Z(new_n1215));
  INV_X1    g1015(.A(G128), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n817), .A2(new_n1216), .B1(new_n249), .B2(new_n815), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(G137), .B2(new_n821), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1159), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n802), .A2(G125), .B1(new_n804), .B2(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1218), .B(new_n1220), .C1(new_n876), .C2(new_n825), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1221), .A2(KEYINPUT59), .ZN(new_n1222));
  AOI211_X1 g1022(.A(G33), .B(G41), .C1(new_n812), .C2(G124), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n829), .B2(new_n354), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1224), .B1(new_n1221), .B2(KEYINPUT59), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1222), .A2(new_n1225), .B1(new_n1211), .B2(new_n1213), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n839), .B1(new_n1215), .B2(new_n1226), .ZN(new_n1227));
  AOI211_X1 g1027(.A(new_n775), .B(new_n1227), .C1(new_n241), .C2(new_n861), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1204), .A2(new_n1228), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT122), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n938), .A2(KEYINPUT40), .B1(new_n950), .B2(new_n951), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1203), .B1(new_n1232), .B2(new_n710), .ZN(new_n1233));
  AND2_X1   g1033(.A1(new_n950), .A2(new_n951), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT40), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1235), .B1(new_n951), .B2(new_n931), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G330), .B(new_n1202), .C1(new_n1234), .C2(new_n1236), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1233), .A2(new_n1237), .A3(new_n970), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n970), .B1(new_n1233), .B2(new_n1237), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1231), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n970), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1202), .B1(new_n953), .B2(G330), .ZN(new_n1242));
  NOR3_X1   g1042(.A1(new_n1232), .A2(new_n710), .A3(new_n1203), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1241), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1233), .A2(new_n1237), .A3(new_n970), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1244), .A2(KEYINPUT122), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1240), .A2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1230), .B1(new_n1247), .B2(new_n1026), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(KEYINPUT57), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1239), .A2(KEYINPUT123), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1251), .B1(new_n1252), .B2(KEYINPUT123), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n716), .B1(new_n1250), .B2(new_n1253), .ZN(new_n1254));
  AOI21_X1  g1054(.A(KEYINPUT57), .B1(new_n1247), .B2(new_n1249), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1248), .B1(new_n1254), .B2(new_n1255), .ZN(G375));
  NAND3_X1  g1056(.A1(new_n1176), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1257));
  NAND3_X1  g1057(.A1(new_n1185), .A2(new_n1046), .A3(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1117), .A2(new_n780), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n271), .B1(new_n812), .B2(G303), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1062), .B(new_n1260), .C1(new_n820), .C2(new_n318), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(G283), .B2(new_n871), .ZN(new_n1262));
  AOI22_X1  g1062(.A1(G116), .A2(new_n807), .B1(new_n802), .B2(G294), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n804), .A2(G97), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1262), .A2(new_n1263), .A3(new_n996), .A4(new_n1264), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n825), .A2(new_n1159), .B1(new_n817), .B2(new_n873), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n1266), .B1(G132), .B2(new_n802), .ZN(new_n1267));
  XOR2_X1   g1067(.A(new_n1267), .B(KEYINPUT124), .Z(new_n1268));
  AOI21_X1  g1068(.A(new_n347), .B1(new_n812), .B2(G128), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n241), .B2(new_n815), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(new_n821), .B2(G150), .ZN(new_n1271));
  OAI221_X1 g1071(.A(new_n1271), .B1(new_n835), .B2(new_n829), .C1(new_n354), .C2(new_n805), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1265), .B1(new_n1268), .B2(new_n1272), .ZN(new_n1273));
  AND2_X1   g1073(.A1(new_n1273), .A2(new_n790), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n775), .B(new_n1274), .C1(new_n243), .C2(new_n861), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1181), .A2(new_n1026), .B1(new_n1259), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1258), .A2(new_n1276), .ZN(G381));
  INV_X1    g1077(.A(new_n1011), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1279), .A2(new_n1112), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1024), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1023), .B(new_n1281), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1278), .B1(new_n1280), .B2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1113), .B1(new_n1043), .B2(new_n1088), .ZN(new_n1284));
  OR2_X1    g1084(.A1(G393), .A2(G396), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1283), .A2(new_n883), .A3(new_n1284), .A4(new_n1286), .ZN(new_n1287));
  AND2_X1   g1087(.A1(new_n1142), .A2(new_n1164), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n1189), .B2(new_n1192), .ZN(new_n1289));
  OR4_X1    g1089(.A1(G375), .A2(new_n1287), .A3(G381), .A4(new_n1289), .ZN(G407));
  NOR3_X1   g1090(.A1(new_n1238), .A2(new_n1239), .A3(new_n1231), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT122), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1292));
  OAI21_X1  g1092(.A(new_n1026), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1229), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT57), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1296), .B1(new_n1191), .B2(new_n1184), .ZN(new_n1298));
  OAI21_X1  g1098(.A(KEYINPUT123), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1299));
  OR2_X1    g1099(.A1(new_n1239), .A2(KEYINPUT123), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1086), .B1(new_n1298), .B2(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1294), .B1(new_n1297), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1289), .ZN(new_n1304));
  INV_X1    g1104(.A(G213), .ZN(new_n1305));
  NOR2_X1   g1105(.A1(new_n1305), .A2(G343), .ZN(new_n1306));
  NAND3_X1  g1106(.A1(new_n1303), .A2(new_n1304), .A3(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(G407), .A2(G213), .A3(new_n1307), .ZN(G409));
  INV_X1    g1108(.A(KEYINPUT125), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT60), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1257), .B1(new_n1190), .B2(new_n1310), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1176), .A2(KEYINPUT60), .A3(new_n1183), .A4(new_n1180), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1311), .A2(new_n716), .A3(new_n1312), .ZN(new_n1313));
  AND3_X1   g1113(.A1(new_n1313), .A2(G384), .A3(new_n1276), .ZN(new_n1314));
  AOI21_X1  g1114(.A(G384), .B1(new_n1313), .B2(new_n1276), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1309), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1313), .A2(new_n1276), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n883), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1313), .A2(G384), .A3(new_n1276), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1318), .A2(KEYINPUT125), .A3(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1306), .A2(G2897), .ZN(new_n1321));
  NAND3_X1  g1121(.A1(new_n1316), .A2(new_n1320), .A3(new_n1321), .ZN(new_n1322));
  NOR2_X1   g1122(.A1(new_n1314), .A2(new_n1315), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1323), .A2(KEYINPUT125), .A3(G2897), .A4(new_n1306), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1247), .A2(new_n1046), .A3(new_n1249), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1230), .B1(new_n1301), .B2(new_n1026), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1289), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1328), .B1(G378), .B2(new_n1303), .ZN(new_n1329));
  OAI21_X1  g1129(.A(new_n1325), .B1(new_n1329), .B2(new_n1306), .ZN(new_n1330));
  INV_X1    g1130(.A(KEYINPUT126), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1306), .ZN(new_n1332));
  AOI21_X1  g1132(.A(G375), .B1(new_n1196), .B2(new_n1194), .ZN(new_n1333));
  OAI211_X1 g1133(.A(new_n1332), .B(new_n1323), .C1(new_n1333), .C2(new_n1328), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  AOI22_X1  g1135(.A1(new_n1330), .A2(new_n1331), .B1(new_n1334), .B2(new_n1335), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT127), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(G393), .A2(G396), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1337), .B1(new_n1285), .B2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  NAND3_X1  g1140(.A1(new_n1285), .A2(new_n1337), .A3(new_n1338), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(G390), .A2(new_n1340), .A3(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1341), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1284), .B1(new_n1343), .B2(new_n1339), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1342), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(G387), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1283), .A2(new_n1342), .A3(new_n1344), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT61), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1346), .A2(new_n1347), .A3(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1323), .ZN(new_n1350));
  NOR3_X1   g1150(.A1(new_n1329), .A2(new_n1306), .A3(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1349), .B1(new_n1351), .B2(KEYINPUT63), .ZN(new_n1352));
  OAI211_X1 g1152(.A(KEYINPUT126), .B(new_n1325), .C1(new_n1329), .C2(new_n1306), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1336), .A2(new_n1352), .A3(new_n1353), .ZN(new_n1354));
  NAND2_X1  g1154(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1196), .ZN(new_n1356));
  OAI21_X1  g1156(.A(new_n716), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1357), .A2(KEYINPUT116), .ZN(new_n1358));
  NAND3_X1  g1158(.A1(new_n1358), .A2(new_n1188), .A3(new_n1187), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1195), .B1(new_n1359), .B2(new_n1167), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1303), .B1(new_n1356), .B2(new_n1360), .ZN(new_n1361));
  INV_X1    g1161(.A(new_n1328), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1361), .A2(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT62), .ZN(new_n1364));
  NAND4_X1  g1164(.A1(new_n1363), .A2(new_n1364), .A3(new_n1332), .A4(new_n1323), .ZN(new_n1365));
  NAND3_X1  g1165(.A1(new_n1365), .A2(new_n1348), .A3(new_n1330), .ZN(new_n1366));
  NOR2_X1   g1166(.A1(new_n1329), .A2(new_n1306), .ZN(new_n1367));
  AOI21_X1  g1167(.A(new_n1364), .B1(new_n1367), .B2(new_n1323), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1355), .B1(new_n1366), .B2(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1354), .A2(new_n1369), .ZN(G405));
  NAND2_X1  g1170(.A1(G375), .A2(new_n1304), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1361), .A2(new_n1371), .ZN(new_n1372));
  XNOR2_X1  g1172(.A(new_n1372), .B(new_n1323), .ZN(new_n1373));
  XNOR2_X1  g1173(.A(new_n1373), .B(new_n1355), .ZN(G402));
endmodule


