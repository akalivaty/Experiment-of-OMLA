//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  XNOR2_X1  g000(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(G101), .ZN(new_n188));
  NOR2_X1   g002(.A1(G237), .A2(G953), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G210), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n188), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  OR2_X1    g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n196), .B1(new_n198), .B2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n193), .A2(new_n195), .A3(new_n199), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT64), .A2(G131), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n206), .A2(new_n209), .A3(new_n207), .A4(new_n211), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n213), .A2(KEYINPUT65), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT65), .B1(new_n213), .B2(new_n214), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n203), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n193), .A3(new_n195), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n192), .A3(G143), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n194), .B(G146), .C1(new_n218), .C2(KEYINPUT1), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT66), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n220), .A2(KEYINPUT66), .A3(new_n221), .A4(new_n222), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n210), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n208), .A2(G134), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n207), .A2(new_n230), .A3(G131), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(G116), .B(G119), .Z(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT2), .B(G113), .ZN(new_n235));
  XOR2_X1   g049(.A(new_n234), .B(new_n235), .Z(new_n236));
  NAND3_X1  g050(.A1(new_n217), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  AND3_X1   g051(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(new_n229), .B2(new_n231), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n213), .A2(new_n214), .B1(new_n201), .B2(new_n202), .ZN(new_n240));
  NOR3_X1   g054(.A1(new_n239), .A2(new_n240), .A3(KEYINPUT30), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n217), .A2(new_n233), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(KEYINPUT30), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n191), .B(new_n237), .C1(new_n243), .C2(new_n236), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n236), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n248), .B1(new_n217), .B2(new_n233), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n247), .B1(new_n249), .B2(new_n241), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n250), .A2(KEYINPUT67), .A3(new_n191), .A4(new_n237), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n246), .A2(KEYINPUT31), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT31), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n244), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n237), .A2(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n217), .A2(new_n233), .A3(KEYINPUT28), .A4(new_n236), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n247), .B1(new_n239), .B2(new_n240), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n191), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G472), .ZN(new_n264));
  INV_X1    g078(.A(G902), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT32), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(G902), .B1(new_n255), .B2(new_n262), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT32), .A3(new_n264), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT68), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n250), .A2(new_n237), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n271), .B1(new_n272), .B2(new_n261), .ZN(new_n273));
  AOI211_X1 g087(.A(KEYINPUT68), .B(new_n191), .C1(new_n250), .C2(new_n237), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n275), .B1(new_n260), .B2(new_n261), .ZN(new_n276));
  NOR3_X1   g090(.A1(new_n273), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n237), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n236), .B1(new_n217), .B2(new_n233), .ZN(new_n279));
  OAI211_X1 g093(.A(KEYINPUT69), .B(KEYINPUT28), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n279), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n256), .B1(new_n281), .B2(new_n237), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n237), .B2(new_n256), .ZN(new_n284));
  OAI211_X1 g098(.A(new_n280), .B(KEYINPUT29), .C1(new_n282), .C2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n265), .B1(new_n285), .B2(new_n261), .ZN(new_n286));
  OAI21_X1  g100(.A(G472), .B1(new_n277), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT70), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT70), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n289), .B(G472), .C1(new_n277), .C2(new_n286), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n268), .A2(new_n270), .A3(new_n288), .A4(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT76), .B(KEYINPUT25), .ZN(new_n292));
  XNOR2_X1  g106(.A(KEYINPUT22), .B(G137), .ZN(new_n293));
  XNOR2_X1  g107(.A(new_n293), .B(KEYINPUT74), .ZN(new_n294));
  INV_X1    g108(.A(G953), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n295), .A2(G221), .A3(G234), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n294), .B(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n298));
  INV_X1    g112(.A(G119), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(G128), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n218), .A2(KEYINPUT23), .A3(G119), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n300), .B(new_n301), .C1(G119), .C2(new_n218), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G110), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT24), .B(G110), .Z(new_n304));
  XNOR2_X1  g118(.A(G119), .B(G128), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n303), .A2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT71), .B(G125), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT16), .ZN(new_n309));
  INV_X1    g123(.A(G140), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G125), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(KEYINPUT71), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT71), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G125), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n316), .A3(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n310), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n309), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n192), .B1(new_n312), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(G125), .A2(G140), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n321), .B1(new_n308), .B2(G140), .ZN(new_n322));
  OAI211_X1 g136(.A(G146), .B(new_n311), .C1(new_n322), .C2(new_n309), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n307), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  OAI22_X1  g138(.A1(new_n302), .A2(G110), .B1(new_n305), .B2(new_n304), .ZN(new_n325));
  NAND2_X1  g139(.A1(G125), .A2(G140), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n318), .A2(KEYINPUT72), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT72), .B1(new_n318), .B2(new_n326), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n192), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n323), .A2(new_n325), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT73), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n323), .A2(new_n333), .A3(new_n325), .A4(new_n330), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n324), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n297), .B1(new_n335), .B2(KEYINPUT75), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT75), .ZN(new_n337));
  AOI211_X1 g151(.A(new_n337), .B(new_n324), .C1(new_n332), .C2(new_n334), .ZN(new_n338));
  NOR2_X1   g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n332), .A2(new_n334), .ZN(new_n340));
  INV_X1    g154(.A(new_n324), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NOR3_X1   g156(.A1(new_n342), .A2(new_n337), .A3(new_n297), .ZN(new_n343));
  OAI211_X1 g157(.A(new_n265), .B(new_n292), .C1(new_n339), .C2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G217), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(G234), .B2(new_n265), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n342), .A2(new_n337), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n335), .A2(KEYINPUT75), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(new_n297), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n336), .A2(new_n338), .ZN(new_n350));
  AOI21_X1  g164(.A(G902), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT76), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT25), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n344), .B(new_n346), .C1(new_n351), .C2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT77), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n353), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n339), .A2(new_n343), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n357), .B1(new_n358), .B2(G902), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n359), .A2(KEYINPUT77), .A3(new_n346), .A4(new_n344), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n346), .A2(G902), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n361), .B(KEYINPUT78), .Z(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n339), .B2(new_n343), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n356), .A2(new_n360), .A3(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT9), .B(G234), .ZN(new_n367));
  OAI21_X1  g181(.A(G221), .B1(new_n367), .B2(G902), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n368), .B(KEYINPUT79), .ZN(new_n369));
  INV_X1    g183(.A(G104), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT3), .B1(new_n370), .B2(G107), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n372));
  INV_X1    g186(.A(G107), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n372), .A2(new_n373), .A3(G104), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(G107), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n371), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT80), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT80), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n371), .A2(new_n374), .A3(new_n378), .A4(new_n375), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n377), .A2(G101), .A3(new_n379), .ZN(new_n380));
  OR2_X1    g194(.A1(new_n376), .A2(G101), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT4), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n377), .A2(new_n383), .A3(G101), .A4(new_n379), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT81), .ZN(new_n385));
  AND2_X1   g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n384), .A2(new_n385), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n203), .B(new_n382), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n215), .A2(new_n216), .ZN(new_n389));
  INV_X1    g203(.A(new_n375), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n370), .A2(G107), .ZN(new_n391));
  OAI21_X1  g205(.A(G101), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n381), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT10), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n395), .B1(new_n225), .B2(new_n226), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n381), .A2(new_n223), .A3(new_n392), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n394), .A2(new_n396), .B1(new_n397), .B2(new_n395), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n388), .A2(new_n389), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n393), .A2(new_n238), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(new_n397), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n213), .A2(new_n214), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT12), .ZN(new_n404));
  INV_X1    g218(.A(new_n389), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT12), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n405), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n404), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(G110), .B(G140), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n295), .A2(G227), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT82), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n388), .A2(new_n398), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n405), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n399), .A3(new_n411), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n413), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n414), .B1(new_n413), .B2(new_n417), .ZN(new_n419));
  OAI21_X1  g233(.A(G469), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G469), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(new_n265), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n388), .A2(new_n389), .A3(new_n398), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n389), .B1(new_n388), .B2(new_n398), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n412), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n399), .A2(new_n411), .A3(new_n404), .A4(new_n407), .ZN(new_n426));
  AOI21_X1  g240(.A(G902), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n422), .B1(new_n427), .B2(new_n421), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n369), .B1(new_n420), .B2(new_n428), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n193), .A2(new_n195), .B1(new_n197), .B2(new_n199), .ZN(new_n430));
  INV_X1    g244(.A(new_n202), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n308), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n314), .A2(new_n316), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n223), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G224), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(G953), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n437), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n439), .B1(new_n432), .B2(new_n434), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n437), .A2(KEYINPUT7), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n438), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n435), .A2(KEYINPUT7), .A3(new_n437), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n247), .B(new_n382), .C1(new_n386), .C2(new_n387), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT5), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n299), .A3(G116), .ZN(new_n447));
  OAI211_X1 g261(.A(G113), .B(new_n447), .C1(new_n234), .C2(new_n446), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n448), .B1(new_n234), .B2(new_n235), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n449), .A2(new_n393), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G110), .B(G122), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n445), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n452), .B(KEYINPUT8), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n449), .A2(new_n393), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n454), .B1(new_n455), .B2(new_n450), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT85), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(KEYINPUT85), .B(new_n454), .C1(new_n455), .C2(new_n450), .ZN(new_n459));
  NAND4_X1  g273(.A1(new_n444), .A2(new_n453), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  AND2_X1   g274(.A1(new_n460), .A2(new_n265), .ZN(new_n461));
  OAI21_X1  g275(.A(G210), .B1(G237), .B2(G902), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT6), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(KEYINPUT84), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n445), .A2(new_n451), .ZN(new_n465));
  INV_X1    g279(.A(new_n452), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n464), .ZN(new_n468));
  AOI211_X1 g282(.A(new_n452), .B(new_n468), .C1(new_n445), .C2(new_n451), .ZN(new_n469));
  INV_X1    g283(.A(new_n453), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  OR2_X1    g285(.A1(new_n438), .A2(new_n440), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n461), .B(new_n462), .C1(new_n471), .C2(new_n472), .ZN(new_n473));
  OR2_X1    g287(.A1(new_n473), .A2(KEYINPUT86), .ZN(new_n474));
  INV_X1    g288(.A(new_n462), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n467), .A2(new_n469), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n472), .B1(new_n476), .B2(new_n453), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n460), .A2(new_n265), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n475), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(KEYINPUT86), .A3(new_n473), .ZN(new_n480));
  OAI21_X1  g294(.A(G214), .B1(G237), .B2(G902), .ZN(new_n481));
  XOR2_X1   g295(.A(new_n481), .B(KEYINPUT83), .Z(new_n482));
  AND4_X1   g296(.A1(new_n429), .A2(new_n474), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G475), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n320), .A2(new_n323), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT89), .ZN(new_n486));
  INV_X1    g300(.A(G237), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n487), .A2(new_n295), .A3(G214), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n194), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n189), .A2(G143), .A3(G214), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n486), .B1(new_n491), .B2(G131), .ZN(new_n492));
  AOI211_X1 g306(.A(KEYINPUT89), .B(new_n228), .C1(new_n489), .C2(new_n490), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT17), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n189), .A2(G143), .A3(G214), .ZN(new_n495));
  AOI21_X1  g309(.A(G143), .B1(new_n189), .B2(G214), .ZN(new_n496));
  OAI21_X1  g310(.A(G131), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(KEYINPUT89), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n491), .A2(new_n486), .A3(G131), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n489), .A2(new_n228), .A3(new_n490), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT88), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n489), .A2(KEYINPUT88), .A3(new_n228), .A4(new_n490), .ZN(new_n503));
  NAND4_X1  g317(.A1(new_n498), .A2(new_n499), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n485), .B(new_n494), .C1(KEYINPUT17), .C2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n329), .ZN(new_n506));
  AOI21_X1  g320(.A(G146), .B1(new_n506), .B2(new_n327), .ZN(new_n507));
  AND3_X1   g321(.A1(new_n317), .A2(G146), .A3(new_n318), .ZN(new_n508));
  AND4_X1   g322(.A1(KEYINPUT18), .A2(new_n489), .A3(G131), .A4(new_n490), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n489), .A2(new_n490), .B1(KEYINPUT18), .B2(G131), .ZN(new_n510));
  OAI22_X1  g324(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT87), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT87), .ZN(new_n513));
  OAI221_X1 g327(.A(new_n513), .B1(new_n509), .B2(new_n510), .C1(new_n507), .C2(new_n508), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(G113), .B(G122), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(new_n370), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n505), .A2(new_n515), .A3(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n492), .A2(new_n493), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n519), .A2(KEYINPUT90), .A3(new_n502), .A4(new_n503), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT90), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n504), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT19), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n328), .B2(new_n329), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n317), .A2(KEYINPUT19), .A3(new_n318), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n192), .A3(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n526), .A2(new_n323), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n520), .A2(new_n522), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n517), .B1(new_n528), .B2(new_n515), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n484), .B(new_n265), .C1(new_n518), .C2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT20), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n528), .A2(new_n515), .ZN(new_n533));
  INV_X1    g347(.A(new_n517), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n505), .A2(new_n515), .A3(new_n517), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n537), .A2(KEYINPUT20), .A3(new_n484), .A4(new_n265), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n517), .B1(new_n505), .B2(new_n515), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n265), .B1(new_n518), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G475), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n532), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(G234), .A2(G237), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n543), .A2(G952), .A3(new_n295), .ZN(new_n544));
  XOR2_X1   g358(.A(new_n544), .B(KEYINPUT94), .Z(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT21), .B(G898), .Z(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(KEYINPUT95), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n543), .A2(G902), .A3(G953), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n546), .B1(new_n549), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT93), .ZN(new_n553));
  XNOR2_X1  g367(.A(G116), .B(G122), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n373), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n554), .A2(new_n373), .ZN(new_n557));
  OAI21_X1  g371(.A(KEYINPUT91), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(G128), .B(G143), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n205), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(KEYINPUT13), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n194), .A2(G128), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n561), .B(G134), .C1(KEYINPUT13), .C2(new_n562), .ZN(new_n563));
  XOR2_X1   g377(.A(G116), .B(G122), .Z(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(G107), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT91), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n555), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n558), .A2(new_n560), .A3(new_n563), .A4(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n559), .B(new_n205), .ZN(new_n569));
  INV_X1    g383(.A(G116), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(KEYINPUT14), .A3(G122), .ZN(new_n571));
  OAI211_X1 g385(.A(G107), .B(new_n571), .C1(new_n564), .C2(KEYINPUT14), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n569), .A2(new_n572), .A3(new_n555), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n367), .A2(new_n345), .A3(G953), .ZN(new_n574));
  AND3_X1   g388(.A1(new_n568), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n574), .B1(new_n568), .B2(new_n573), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n553), .B(new_n265), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT92), .ZN(new_n578));
  INV_X1    g392(.A(G478), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n579), .A2(KEYINPUT15), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n568), .A2(new_n573), .ZN(new_n581));
  INV_X1    g395(.A(new_n574), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n568), .A2(new_n573), .A3(new_n574), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT92), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n586), .A3(new_n265), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n578), .A2(new_n580), .A3(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n577), .B(KEYINPUT92), .C1(KEYINPUT15), .C2(new_n579), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n542), .A2(new_n552), .A3(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n291), .A2(new_n366), .A3(new_n483), .A4(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(G101), .ZN(G3));
  AOI22_X1  g407(.A1(new_n252), .A2(new_n254), .B1(new_n261), .B2(new_n260), .ZN(new_n594));
  OAI21_X1  g408(.A(G472), .B1(new_n594), .B2(G902), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n266), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n369), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n413), .A2(new_n417), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n598), .A2(KEYINPUT82), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n413), .A2(new_n414), .A3(new_n417), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n421), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n427), .A2(new_n421), .ZN(new_n602));
  INV_X1    g416(.A(new_n422), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n597), .B1(new_n601), .B2(new_n604), .ZN(new_n605));
  NOR3_X1   g419(.A1(new_n596), .A2(new_n365), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n479), .A2(new_n473), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n481), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT97), .B(G478), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n575), .A2(new_n576), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(G902), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n612));
  OAI21_X1  g426(.A(KEYINPUT33), .B1(new_n576), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n610), .A2(new_n613), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n265), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n611), .B1(new_n617), .B2(new_n579), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n542), .A2(new_n618), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n608), .A2(new_n552), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n606), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT34), .B(G104), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(KEYINPUT98), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n621), .B(new_n623), .ZN(G6));
  NAND4_X1  g438(.A1(new_n590), .A2(new_n541), .A3(new_n532), .A4(new_n538), .ZN(new_n625));
  XOR2_X1   g439(.A(new_n552), .B(KEYINPUT99), .Z(new_n626));
  NOR3_X1   g440(.A1(new_n608), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n606), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  INV_X1    g444(.A(new_n596), .ZN(new_n631));
  INV_X1    g445(.A(new_n297), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n632), .A2(KEYINPUT36), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n342), .B(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(new_n363), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n356), .A2(new_n360), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n483), .A2(new_n591), .A3(new_n631), .A4(new_n636), .ZN(new_n637));
  XOR2_X1   g451(.A(new_n637), .B(KEYINPUT37), .Z(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G110), .ZN(G12));
  INV_X1    g453(.A(new_n481), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n640), .B1(new_n479), .B2(new_n473), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n545), .B1(G900), .B2(new_n550), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n625), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g458(.A1(new_n429), .A2(new_n641), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n291), .A2(new_n636), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G128), .ZN(G30));
  AND2_X1   g461(.A1(new_n246), .A2(new_n251), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n281), .A2(new_n237), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n648), .B1(new_n261), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(G472), .B1(new_n650), .B2(G902), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n268), .A2(new_n270), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(KEYINPUT100), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT32), .B1(new_n269), .B2(new_n264), .ZN(new_n654));
  NOR4_X1   g468(.A1(new_n594), .A2(new_n267), .A3(G472), .A4(G902), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT100), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n656), .A2(new_n657), .A3(new_n651), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n356), .A2(new_n360), .A3(new_n635), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n481), .ZN(new_n661));
  XOR2_X1   g475(.A(new_n642), .B(KEYINPUT39), .Z(new_n662));
  NOR2_X1   g476(.A1(new_n605), .A2(new_n662), .ZN(new_n663));
  OR2_X1    g477(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n542), .A2(new_n590), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n480), .A2(new_n474), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT38), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n659), .A2(new_n666), .A3(new_n668), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G143), .ZN(G45));
  NOR2_X1   g487(.A1(new_n608), .A2(new_n605), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n619), .A2(new_n643), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n291), .A2(new_n636), .A3(new_n674), .A4(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G146), .ZN(G48));
  INV_X1    g491(.A(new_n602), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n427), .A2(new_n421), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n597), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n291), .A2(new_n620), .A3(new_n366), .A4(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(KEYINPUT41), .B(G113), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G15));
  NAND4_X1  g499(.A1(new_n291), .A2(new_n627), .A3(new_n366), .A4(new_n682), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G116), .ZN(G18));
  NOR2_X1   g501(.A1(new_n681), .A2(new_n608), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n291), .A2(new_n591), .A3(new_n636), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  OAI21_X1  g504(.A(new_n280), .B1(new_n282), .B2(new_n284), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n261), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n255), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n693), .A2(KEYINPUT101), .A3(new_n264), .A4(new_n265), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT101), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n252), .A2(new_n254), .B1(new_n691), .B2(new_n261), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n264), .A2(new_n265), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n695), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n694), .A2(new_n595), .A3(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(new_n626), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n641), .A2(new_n700), .A3(new_n668), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n699), .A2(new_n701), .A3(new_n366), .A4(new_n682), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT102), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G122), .ZN(G24));
  NAND4_X1  g518(.A1(new_n699), .A2(new_n688), .A3(new_n636), .A4(new_n675), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT103), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n313), .ZN(G27));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n708));
  AOI211_X1 g522(.A(new_n369), .B(new_n640), .C1(new_n480), .C2(new_n474), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n598), .A2(KEYINPUT104), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT104), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n417), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n710), .A2(G469), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n428), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n291), .A2(new_n709), .A3(new_n366), .A4(new_n714), .ZN(new_n715));
  INV_X1    g529(.A(new_n675), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n708), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n654), .B1(KEYINPUT105), .B2(new_n270), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n288), .A2(new_n290), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  OR2_X1    g534(.A1(new_n270), .A2(KEYINPUT105), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n669), .A2(new_n597), .A3(new_n481), .A4(new_n714), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n723), .A2(new_n716), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n722), .A2(new_n724), .A3(KEYINPUT42), .A4(new_n366), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n717), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G131), .ZN(G33));
  NOR3_X1   g541(.A1(new_n719), .A2(new_n654), .A3(new_n655), .ZN(new_n728));
  INV_X1    g542(.A(new_n644), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n728), .A2(new_n723), .A3(new_n365), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(new_n205), .ZN(G36));
  NAND2_X1  g545(.A1(new_n669), .A2(new_n481), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n618), .A2(new_n541), .A3(new_n532), .A4(new_n538), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n734), .B(KEYINPUT43), .Z(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n596), .A3(new_n636), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n733), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n599), .A2(new_n600), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n741), .A2(KEYINPUT45), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n710), .A2(KEYINPUT45), .A3(new_n712), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n742), .A2(new_n743), .A3(KEYINPUT106), .A4(G469), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n743), .B(G469), .C1(new_n741), .C2(KEYINPUT45), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n422), .B1(new_n744), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n602), .B1(new_n748), .B2(KEYINPUT46), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT46), .ZN(new_n750));
  AOI211_X1 g564(.A(new_n750), .B(new_n422), .C1(new_n744), .C2(new_n747), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n597), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n662), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n736), .A2(new_n737), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n740), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G137), .ZN(G39));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  OAI211_X1 g572(.A(KEYINPUT47), .B(new_n597), .C1(new_n749), .C2(new_n751), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n291), .A2(new_n366), .A3(new_n716), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n733), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G140), .ZN(G42));
  INV_X1    g577(.A(KEYINPUT52), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n676), .A2(new_n646), .A3(new_n705), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n652), .A2(new_n597), .A3(new_n660), .A4(new_n642), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n641), .A2(new_n668), .A3(new_n714), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n764), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n660), .B1(new_n656), .B2(new_n720), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n694), .A2(new_n595), .A3(new_n698), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n771), .A2(new_n660), .A3(new_n716), .ZN(new_n772));
  AOI22_X1  g586(.A1(new_n770), .A2(new_n645), .B1(new_n772), .B2(new_n688), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n636), .B1(new_n656), .B2(new_n651), .ZN(new_n774));
  INV_X1    g588(.A(new_n767), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n774), .A2(new_n597), .A3(new_n642), .A4(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n773), .A2(KEYINPUT52), .A3(new_n776), .A4(new_n676), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n769), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT53), .B1(new_n778), .B2(KEYINPUT109), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n683), .A2(new_n686), .A3(new_n689), .A4(new_n702), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n420), .A2(new_n428), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n542), .A2(new_n590), .A3(new_n643), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n291), .A2(new_n709), .A3(new_n781), .A4(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n709), .A2(new_n699), .A3(new_n675), .A4(new_n714), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n780), .B1(new_n636), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n619), .A2(new_n625), .ZN(new_n787));
  AND4_X1   g601(.A1(new_n474), .A2(new_n787), .A3(new_n480), .A4(new_n482), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n365), .A2(new_n605), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n788), .A2(new_n631), .A3(new_n789), .A4(new_n700), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n592), .A2(new_n637), .A3(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n730), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n778), .A2(new_n726), .A3(new_n786), .A4(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n779), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT54), .ZN(new_n795));
  XNOR2_X1  g609(.A(KEYINPUT110), .B(KEYINPUT54), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n769), .A2(new_n777), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n785), .A2(new_n636), .ZN(new_n798));
  AND4_X1   g612(.A1(new_n683), .A2(new_n686), .A3(new_n689), .A4(new_n702), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n726), .A2(new_n792), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  OAI21_X1  g614(.A(KEYINPUT53), .B1(new_n797), .B2(new_n800), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n726), .A2(new_n792), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n802), .A2(new_n778), .A3(new_n803), .A4(new_n786), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n796), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n735), .A2(new_n546), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n699), .A2(new_n366), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  XNOR2_X1  g623(.A(new_n680), .B(KEYINPUT111), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n810), .A2(new_n369), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n733), .B(new_n809), .C1(new_n760), .C2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n808), .A2(new_n681), .ZN(new_n813));
  AND2_X1   g627(.A1(new_n735), .A2(new_n546), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT50), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n481), .B1(KEYINPUT112), .B2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n813), .A2(new_n814), .A3(new_n670), .A4(new_n816), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n815), .A2(KEYINPUT112), .ZN(new_n818));
  INV_X1    g632(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n807), .A2(new_n808), .A3(new_n681), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n670), .A3(new_n818), .A4(new_n816), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n732), .A2(new_n545), .A3(new_n681), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n735), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n699), .A2(new_n636), .ZN(new_n826));
  OR3_X1    g640(.A1(new_n825), .A2(KEYINPUT113), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT113), .B1(new_n825), .B2(new_n826), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n659), .A2(new_n365), .ZN(new_n830));
  INV_X1    g644(.A(new_n542), .ZN(new_n831));
  INV_X1    g645(.A(new_n618), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n824), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n823), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n812), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(KEYINPUT51), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n812), .A2(new_n834), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n722), .A2(new_n366), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n825), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n841), .B(KEYINPUT48), .Z(new_n842));
  NAND4_X1  g656(.A1(new_n830), .A2(new_n542), .A3(new_n618), .A4(new_n824), .ZN(new_n843));
  INV_X1    g657(.A(G952), .ZN(new_n844));
  AOI211_X1 g658(.A(new_n844), .B(G953), .C1(new_n809), .C2(new_n688), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n842), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n795), .A2(new_n806), .A3(new_n839), .A4(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT114), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n844), .A2(new_n295), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n805), .B1(new_n794), .B2(KEYINPUT54), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(KEYINPUT114), .A3(new_n846), .A4(new_n839), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n849), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n482), .ZN(new_n854));
  INV_X1    g668(.A(new_n680), .ZN(new_n855));
  AOI211_X1 g669(.A(new_n854), .B(new_n671), .C1(KEYINPUT49), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(KEYINPUT49), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT108), .Z(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n365), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n659), .A2(new_n734), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n856), .A2(new_n597), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n853), .A2(new_n861), .ZN(G75));
  INV_X1    g676(.A(KEYINPUT117), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n801), .A2(G902), .A3(new_n804), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT116), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n801), .A2(new_n804), .A3(new_n866), .A4(G902), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n865), .A2(new_n475), .A3(new_n867), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n471), .B(new_n472), .Z(new_n869));
  XOR2_X1   g683(.A(new_n869), .B(KEYINPUT55), .Z(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(KEYINPUT56), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n295), .A2(G952), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n872), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n870), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n801), .A2(new_n804), .A3(G210), .A4(G902), .ZN(new_n877));
  OR2_X1    g691(.A1(new_n877), .A2(KEYINPUT115), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT56), .B1(new_n877), .B2(KEYINPUT115), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n863), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n878), .A2(new_n879), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(new_n870), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n883), .A2(KEYINPUT117), .A3(new_n872), .A4(new_n874), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n881), .A2(new_n884), .ZN(G51));
  AND3_X1   g699(.A1(new_n801), .A2(new_n804), .A3(new_n796), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n886), .A2(new_n805), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT118), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n422), .B(KEYINPUT57), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n425), .A2(new_n426), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n889), .B1(new_n886), .B2(new_n805), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(KEYINPUT118), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n865), .A2(new_n747), .A3(new_n744), .A4(new_n867), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n873), .B1(new_n894), .B2(new_n895), .ZN(G54));
  NAND4_X1  g710(.A1(new_n865), .A2(KEYINPUT58), .A3(G475), .A4(new_n867), .ZN(new_n897));
  INV_X1    g711(.A(new_n537), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n874), .ZN(new_n900));
  OR3_X1    g714(.A1(new_n897), .A2(KEYINPUT119), .A3(new_n898), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT119), .B1(new_n897), .B2(new_n898), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(G60));
  NOR2_X1   g717(.A1(new_n615), .A2(new_n616), .ZN(new_n904));
  NAND2_X1  g718(.A1(G478), .A2(G902), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT59), .Z(new_n906));
  NOR2_X1   g720(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n795), .A2(new_n806), .ZN(new_n908));
  INV_X1    g722(.A(new_n906), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AOI221_X4 g724(.A(new_n873), .B1(new_n887), .B2(new_n907), .C1(new_n910), .C2(new_n904), .ZN(G63));
  NAND2_X1  g725(.A1(new_n801), .A2(new_n804), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT60), .Z(new_n915));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n358), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n913), .A2(new_n634), .A3(new_n915), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n917), .A2(new_n874), .A3(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT120), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT61), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n919), .B(new_n921), .ZN(G66));
  OR2_X1    g736(.A1(new_n780), .A2(new_n791), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n295), .ZN(new_n924));
  OAI21_X1  g738(.A(G953), .B1(new_n549), .B2(new_n436), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT121), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n471), .B1(G898), .B2(new_n295), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n927), .B(new_n928), .Z(G69));
  AND2_X1   g743(.A1(new_n524), .A2(new_n525), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n243), .B(new_n930), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(G900), .A2(G953), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n840), .A2(new_n608), .A3(new_n667), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n765), .B1(new_n753), .B2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n730), .B1(new_n717), .B2(new_n725), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n762), .A2(new_n755), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  OAI211_X1 g751(.A(new_n932), .B(new_n933), .C1(new_n937), .C2(G953), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT122), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT62), .ZN(new_n940));
  INV_X1    g754(.A(new_n672), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(new_n941), .B2(new_n765), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n672), .A2(KEYINPUT62), .A3(new_n676), .A4(new_n773), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n728), .A2(new_n365), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n945), .A2(new_n663), .A3(new_n733), .A4(new_n787), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n944), .A2(new_n762), .A3(new_n755), .A4(new_n946), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n295), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n939), .B1(new_n948), .B2(new_n931), .ZN(new_n949));
  AOI211_X1 g763(.A(KEYINPUT122), .B(new_n932), .C1(new_n947), .C2(new_n295), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n938), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n295), .B1(G227), .B2(G900), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n952), .B1(new_n938), .B2(KEYINPUT123), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  OAI221_X1 g768(.A(new_n938), .B1(KEYINPUT123), .B2(new_n952), .C1(new_n949), .C2(new_n950), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n954), .A2(new_n955), .ZN(G72));
  NAND2_X1  g770(.A1(G472), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT63), .Z(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT124), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n947), .B2(new_n923), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT125), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI211_X1 g776(.A(KEYINPUT125), .B(new_n959), .C1(new_n947), .C2(new_n923), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n962), .A2(new_n191), .A3(new_n272), .A4(new_n963), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n959), .B1(new_n937), .B2(new_n923), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n965), .A2(new_n261), .A3(new_n237), .A4(new_n250), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n964), .A2(new_n874), .A3(new_n966), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n273), .A2(new_n274), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n958), .B1(new_n968), .B2(new_n648), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT126), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n794), .A2(new_n970), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT127), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n967), .A2(new_n972), .ZN(G57));
endmodule


