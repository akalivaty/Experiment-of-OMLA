//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n542, new_n543, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n560, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n571, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n605, new_n606,
    new_n607, new_n608, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n623,
    new_n626, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n839, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1205, new_n1206, new_n1207, new_n1208;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT65), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n462), .B1(new_n463), .B2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n465), .A2(KEYINPUT67), .A3(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(G137), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n463), .A2(G2104), .ZN(new_n469));
  NAND4_X1  g044(.A1(new_n464), .A2(new_n466), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n465), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n470), .A2(KEYINPUT68), .A3(new_n472), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G125), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n463), .A2(G2104), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n480));
  OAI21_X1  g055(.A(KEYINPUT66), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n482));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n482), .A2(new_n469), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n478), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g060(.A1(G113), .A2(G2104), .ZN(new_n486));
  OAI21_X1  g061(.A(G2105), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n477), .A2(new_n487), .ZN(G160));
  NAND3_X1  g063(.A1(new_n464), .A2(new_n469), .A3(new_n466), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT69), .ZN(new_n490));
  XNOR2_X1  g065(.A(new_n489), .B(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G136), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n491), .A2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G124), .ZN(new_n498));
  OR2_X1    g073(.A1(G100), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G112), .C2(new_n492), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n495), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G162));
  INV_X1    g077(.A(G138), .ZN(new_n503));
  NOR3_X1   g078(.A1(new_n503), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n504));
  AND3_X1   g079(.A1(new_n482), .A2(new_n469), .A3(new_n483), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n483), .B1(new_n482), .B2(new_n469), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n503), .A2(G2105), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n464), .A2(new_n466), .A3(new_n508), .A4(new_n469), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT4), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(new_n466), .A2(new_n469), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  AND2_X1   g088(.A1(G126), .A2(G2105), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n512), .A2(new_n513), .A3(new_n464), .A4(new_n514), .ZN(new_n515));
  NAND4_X1  g090(.A1(new_n464), .A2(new_n466), .A3(new_n469), .A4(new_n514), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT70), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g093(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n519));
  INV_X1    g094(.A(G114), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n519), .B1(new_n520), .B2(G2105), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n511), .A2(new_n518), .A3(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(new_n523), .ZN(G164));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  XOR2_X1   g101(.A(new_n526), .B(KEYINPUT71), .Z(new_n527));
  XNOR2_X1  g102(.A(KEYINPUT5), .B(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G62), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n525), .B1(new_n527), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G543), .ZN(new_n531));
  OR2_X1    g106(.A1(KEYINPUT6), .A2(G651), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT6), .A2(G651), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n531), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G50), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n532), .A2(new_n533), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(new_n528), .ZN(new_n537));
  INV_X1    g112(.A(G88), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n535), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n530), .A2(new_n539), .ZN(G303));
  INV_X1    g115(.A(G303), .ZN(G166));
  XNOR2_X1  g116(.A(KEYINPUT72), .B(KEYINPUT7), .ZN(new_n542));
  NAND3_X1  g117(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n542), .B(new_n543), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n536), .A2(new_n528), .ZN(new_n545));
  XNOR2_X1  g120(.A(KEYINPUT73), .B(G89), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(KEYINPUT74), .ZN(new_n548));
  AND2_X1   g123(.A1(G63), .A2(G651), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n534), .A2(G51), .B1(new_n528), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n547), .A2(KEYINPUT74), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(G168));
  NAND2_X1  g128(.A1(new_n534), .A2(G52), .ZN(new_n554));
  INV_X1    g129(.A(G90), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n537), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n528), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n525), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n556), .A2(new_n558), .ZN(G171));
  NAND2_X1  g134(.A1(new_n534), .A2(G43), .ZN(new_n560));
  INV_X1    g135(.A(G81), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n560), .B1(new_n537), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n528), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n563), .A2(new_n525), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G860), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT75), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g143(.A(KEYINPUT76), .B(KEYINPUT8), .Z(new_n569));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n569), .B(new_n570), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  AOI22_X1  g147(.A1(new_n528), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G91), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n573), .A2(new_n525), .B1(new_n537), .B2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT9), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n534), .A2(new_n576), .A3(G53), .ZN(new_n577));
  AND2_X1   g152(.A1(KEYINPUT6), .A2(G651), .ZN(new_n578));
  NOR2_X1   g153(.A1(KEYINPUT6), .A2(G651), .ZN(new_n579));
  OAI211_X1 g154(.A(G53), .B(G543), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n580), .A2(KEYINPUT9), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n577), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n577), .A2(new_n581), .A3(KEYINPUT77), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n575), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(G299));
  INV_X1    g162(.A(G171), .ZN(G301));
  INV_X1    g163(.A(G168), .ZN(G286));
  INV_X1    g164(.A(KEYINPUT78), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n545), .A2(new_n590), .A3(G87), .ZN(new_n591));
  INV_X1    g166(.A(G87), .ZN(new_n592));
  OAI21_X1  g167(.A(KEYINPUT78), .B1(new_n537), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n528), .A2(G74), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G49), .B2(new_n534), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n594), .A2(new_n596), .ZN(G288));
  NAND2_X1  g172(.A1(new_n534), .A2(G48), .ZN(new_n598));
  INV_X1    g173(.A(G86), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n537), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n528), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(new_n525), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(G305));
  XNOR2_X1  g179(.A(KEYINPUT79), .B(G47), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n545), .A2(G85), .B1(new_n534), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT80), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n528), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n525), .B2(new_n608), .ZN(G290));
  NAND2_X1  g184(.A1(G301), .A2(G868), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n545), .A2(G92), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT10), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n612), .B1(G54), .B2(new_n534), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n528), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n614), .A2(KEYINPUT81), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(KEYINPUT81), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n615), .A2(G651), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n610), .B1(new_n619), .B2(G868), .ZN(G284));
  OAI21_X1  g195(.A(new_n610), .B1(new_n619), .B2(G868), .ZN(G321));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(G299), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G168), .B2(new_n622), .ZN(G297));
  OAI21_X1  g199(.A(new_n623), .B1(G168), .B2(new_n622), .ZN(G280));
  INV_X1    g200(.A(G559), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n619), .B1(new_n626), .B2(G860), .ZN(G148));
  NAND2_X1  g202(.A1(new_n619), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G868), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(G868), .B2(new_n565), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n632), .B(G2104), .C1(G111), .C2(new_n492), .ZN(new_n633));
  INV_X1    g208(.A(G135), .ZN(new_n634));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n633), .B1(new_n493), .B2(new_n634), .C1(new_n635), .C2(new_n496), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  OAI21_X1  g212(.A(new_n471), .B1(new_n505), .B2(new_n506), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT12), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2100), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n637), .A2(new_n641), .ZN(G156));
  XOR2_X1   g217(.A(KEYINPUT15), .B(G2435), .Z(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT83), .B(G2438), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2427), .B(G2430), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(KEYINPUT82), .B(KEYINPUT14), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n645), .A2(new_n647), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n648), .A2(new_n649), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2451), .B(G2454), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n651), .B(new_n655), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2443), .B(G2446), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(G14), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n660), .B1(new_n659), .B2(new_n657), .ZN(G401));
  XNOR2_X1  g236(.A(G2067), .B(G2678), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT84), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT85), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n666), .B1(new_n665), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2084), .B(G2090), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n664), .B(KEYINPUT17), .Z(new_n669));
  INV_X1    g244(.A(new_n662), .ZN(new_n670));
  OAI211_X1 g245(.A(new_n667), .B(new_n668), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n670), .A2(new_n668), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n664), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT18), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n662), .A2(new_n668), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n669), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n671), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2096), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G227));
  XOR2_X1   g255(.A(G1971), .B(G1976), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT19), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n682), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n682), .B2(new_n688), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(G229));
  OAI21_X1  g273(.A(KEYINPUT94), .B1(G29), .B2(G32), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n494), .A2(G141), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n497), .A2(G129), .ZN(new_n701));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  INV_X1    g277(.A(KEYINPUT26), .ZN(new_n703));
  OR2_X1    g278(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n702), .A2(new_n703), .ZN(new_n705));
  AOI22_X1  g280(.A1(new_n704), .A2(new_n705), .B1(G105), .B2(new_n471), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n700), .A2(new_n701), .A3(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G29), .ZN(new_n709));
  MUX2_X1   g284(.A(KEYINPUT94), .B(new_n699), .S(new_n709), .Z(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT27), .B(G1996), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G29), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n713), .A2(G33), .ZN(new_n714));
  OAI21_X1  g289(.A(G127), .B1(new_n505), .B2(new_n506), .ZN(new_n715));
  INV_X1    g290(.A(G115), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n465), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n717), .A2(G2105), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n492), .A2(G103), .A3(G2104), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT25), .Z(new_n720));
  INV_X1    g295(.A(G139), .ZN(new_n721));
  OAI211_X1 g296(.A(new_n718), .B(new_n720), .C1(new_n721), .C2(new_n493), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n714), .B1(new_n722), .B2(G29), .ZN(new_n723));
  INV_X1    g298(.A(G2072), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT92), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n712), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G21), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G168), .B2(new_n728), .ZN(new_n730));
  INV_X1    g305(.A(G1966), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n636), .A2(new_n713), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n728), .A2(G5), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G171), .B2(new_n728), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G1961), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT30), .B(G28), .ZN(new_n737));
  OR2_X1    g312(.A1(KEYINPUT31), .A2(G11), .ZN(new_n738));
  NAND2_X1  g313(.A1(KEYINPUT31), .A2(G11), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n737), .A2(new_n713), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND4_X1  g315(.A1(new_n732), .A2(new_n733), .A3(new_n736), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(G164), .A2(G29), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G27), .B2(G29), .ZN(new_n743));
  INV_X1    g318(.A(G2078), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n723), .B2(new_n724), .ZN(new_n746));
  NAND2_X1  g321(.A1(G160), .A2(G29), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT93), .B(KEYINPUT24), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(G34), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n747), .B1(G29), .B2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G2084), .ZN(new_n751));
  OAI22_X1  g326(.A1(new_n750), .A2(new_n751), .B1(new_n743), .B2(new_n744), .ZN(new_n752));
  NOR4_X1   g327(.A1(new_n727), .A2(new_n741), .A3(new_n746), .A4(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n710), .A2(new_n711), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n750), .A2(new_n751), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT95), .Z(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G1961), .B2(new_n735), .ZN(new_n757));
  OAI21_X1  g332(.A(KEYINPUT96), .B1(new_n754), .B2(new_n757), .ZN(new_n758));
  OR3_X1    g333(.A1(new_n754), .A2(new_n757), .A3(KEYINPUT96), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n753), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(KEYINPUT97), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT97), .ZN(new_n762));
  NAND4_X1  g337(.A1(new_n753), .A2(new_n762), .A3(new_n758), .A4(new_n759), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n728), .A2(G19), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(new_n565), .B2(new_n728), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(G1341), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n619), .A2(G16), .ZN(new_n767));
  OAI21_X1  g342(.A(new_n767), .B1(G4), .B2(G16), .ZN(new_n768));
  INV_X1    g343(.A(G1348), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n769), .B2(new_n768), .ZN(new_n771));
  NOR2_X1   g346(.A1(G29), .A2(G35), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G162), .B2(G29), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n773), .B(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G2090), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n728), .A2(G20), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT23), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n586), .B2(new_n728), .ZN(new_n780));
  INV_X1    g355(.A(G1956), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n771), .A2(new_n777), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n713), .A2(G26), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT28), .Z(new_n785));
  OR2_X1    g360(.A1(G104), .A2(G2105), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n786), .B(G2104), .C1(G116), .C2(new_n492), .ZN(new_n787));
  INV_X1    g362(.A(G140), .ZN(new_n788));
  INV_X1    g363(.A(G128), .ZN(new_n789));
  OAI221_X1 g364(.A(new_n787), .B1(new_n493), .B2(new_n788), .C1(new_n789), .C2(new_n496), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT91), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n785), .B1(new_n791), .B2(G29), .ZN(new_n792));
  INV_X1    g367(.A(G2067), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n775), .A2(new_n776), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n783), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n761), .A2(new_n763), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n728), .A2(G22), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G166), .B2(new_n728), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT88), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(G1971), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(G1971), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n728), .A2(G23), .ZN(new_n803));
  AND2_X1   g378(.A1(new_n594), .A2(new_n596), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n803), .B1(new_n804), .B2(new_n728), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT33), .B(G1976), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n728), .A2(G6), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n808), .B1(new_n603), .B2(new_n728), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT32), .B(G1981), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT87), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n809), .B(new_n811), .ZN(new_n812));
  NAND4_X1  g387(.A1(new_n801), .A2(new_n802), .A3(new_n807), .A4(new_n812), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n814));
  MUX2_X1   g389(.A(G24), .B(G290), .S(G16), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G1986), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n813), .B2(KEYINPUT34), .ZN(new_n817));
  OAI21_X1  g392(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n818));
  INV_X1    g393(.A(G107), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n818), .B1(new_n819), .B2(G2105), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(new_n494), .B2(G131), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT86), .ZN(new_n822));
  AND3_X1   g397(.A1(new_n497), .A2(new_n822), .A3(G119), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n822), .B1(new_n497), .B2(G119), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G29), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(G25), .B2(G29), .ZN(new_n828));
  XOR2_X1   g403(.A(KEYINPUT35), .B(G1991), .Z(new_n829));
  OR2_X1    g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n814), .A2(new_n817), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n832), .A2(KEYINPUT36), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT90), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n832), .A2(KEYINPUT36), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT89), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n797), .B1(new_n835), .B2(new_n837), .ZN(G311));
  NAND2_X1  g413(.A1(new_n835), .A2(new_n837), .ZN(new_n839));
  INV_X1    g414(.A(new_n797), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(G150));
  NAND2_X1  g416(.A1(new_n619), .A2(G559), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT38), .ZN(new_n843));
  INV_X1    g418(.A(new_n565), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n534), .A2(G55), .ZN(new_n845));
  INV_X1    g420(.A(G93), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(new_n537), .B2(new_n846), .ZN(new_n847));
  AOI22_X1  g422(.A1(new_n528), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n848), .A2(new_n525), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n844), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n565), .A2(new_n850), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n843), .B(new_n855), .ZN(new_n856));
  OR2_X1    g431(.A1(new_n856), .A2(KEYINPUT39), .ZN(new_n857));
  INV_X1    g432(.A(G860), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(KEYINPUT39), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n850), .A2(new_n858), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT37), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(G145));
  XNOR2_X1  g438(.A(new_n501), .B(G160), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(new_n636), .Z(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT99), .ZN(new_n867));
  INV_X1    g442(.A(new_n722), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n791), .A2(new_n707), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n790), .A2(KEYINPUT91), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n790), .A2(KEYINPUT91), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n708), .A3(new_n871), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n869), .A2(G164), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(G164), .B1(new_n869), .B2(new_n872), .ZN(new_n874));
  OAI211_X1 g449(.A(new_n867), .B(new_n868), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n869), .A2(new_n872), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n523), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n868), .A2(new_n867), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n722), .A2(KEYINPUT99), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n869), .A2(G164), .A3(new_n872), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n877), .A2(new_n878), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n825), .B(new_n639), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n494), .A2(G142), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n497), .A2(G130), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n492), .A2(G118), .ZN(new_n885));
  OAI21_X1  g460(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n883), .B(new_n884), .C1(new_n885), .C2(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n882), .B(new_n887), .Z(new_n888));
  AND3_X1   g463(.A1(new_n875), .A2(new_n881), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n888), .B1(new_n875), .B2(new_n881), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n866), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n875), .A2(new_n881), .ZN(new_n892));
  INV_X1    g467(.A(new_n888), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n875), .A2(new_n881), .A3(new_n888), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n894), .A2(new_n865), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(G37), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n891), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  XOR2_X1   g473(.A(KEYINPUT100), .B(KEYINPUT40), .Z(new_n899));
  XNOR2_X1  g474(.A(new_n898), .B(new_n899), .ZN(G395));
  XNOR2_X1  g475(.A(G288), .B(KEYINPUT101), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n603), .ZN(new_n902));
  XNOR2_X1  g477(.A(G290), .B(G166), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT42), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n904), .A2(KEYINPUT102), .A3(new_n905), .ZN(new_n906));
  XOR2_X1   g481(.A(new_n902), .B(new_n903), .Z(new_n907));
  NOR2_X1   g482(.A1(new_n905), .A2(KEYINPUT102), .ZN(new_n908));
  AND2_X1   g483(.A1(new_n905), .A2(KEYINPUT102), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n618), .A2(G299), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n618), .A2(G299), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT41), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n915), .B1(new_n912), .B2(new_n913), .ZN(new_n916));
  INV_X1    g491(.A(new_n913), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n917), .A2(KEYINPUT41), .A3(new_n911), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n628), .B(new_n855), .ZN(new_n921));
  MUX2_X1   g496(.A(new_n914), .B(new_n920), .S(new_n921), .Z(new_n922));
  AOI211_X1 g497(.A(new_n906), .B(new_n910), .C1(new_n922), .C2(KEYINPUT103), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(KEYINPUT103), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  OAI21_X1  g501(.A(G868), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n851), .A2(new_n622), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n927), .A2(new_n928), .ZN(G295));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n928), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n931));
  XNOR2_X1  g506(.A(G171), .B(KEYINPUT104), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n855), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(new_n932), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n854), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n933), .A2(new_n935), .A3(G168), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n855), .A2(new_n932), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n934), .A2(new_n854), .ZN(new_n938));
  OAI21_X1  g513(.A(G286), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n914), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(new_n936), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n940), .B1(new_n919), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(new_n907), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n904), .B(new_n940), .C1(new_n919), .C2(new_n941), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n943), .A2(new_n944), .A3(new_n897), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT43), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT105), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n931), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT43), .ZN(new_n949));
  NAND4_X1  g524(.A1(new_n943), .A2(new_n944), .A3(new_n949), .A4(new_n897), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  XOR2_X1   g526(.A(new_n948), .B(new_n951), .Z(G397));
  NAND2_X1  g527(.A1(new_n791), .A2(G2067), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n870), .A2(new_n793), .A3(new_n871), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n708), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n521), .B1(new_n507), .B2(new_n510), .ZN(new_n956));
  AOI21_X1  g531(.A(G1384), .B1(new_n956), .B2(new_n518), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n477), .A2(new_n487), .A3(G40), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n957), .A2(new_n958), .A3(KEYINPUT45), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n955), .A2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1996), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n962), .B(KEYINPUT46), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n960), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT125), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT125), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n960), .A2(new_n966), .A3(new_n963), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n965), .A2(KEYINPUT47), .A3(new_n967), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n707), .B(new_n961), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n953), .A2(new_n954), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n826), .A2(new_n829), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n954), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  XOR2_X1   g550(.A(new_n825), .B(new_n829), .Z(new_n976));
  OAI21_X1  g551(.A(new_n959), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g552(.A1(G290), .A2(G1986), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n959), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT48), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n959), .A2(new_n975), .B1(new_n977), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n970), .A2(new_n971), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT126), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT126), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n970), .A2(new_n981), .A3(new_n984), .A4(new_n971), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n477), .A2(new_n487), .A3(G40), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT45), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(G1384), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n523), .A2(new_n989), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n987), .B(new_n990), .C1(KEYINPUT45), .C2(new_n957), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n991), .A2(new_n731), .ZN(new_n992));
  INV_X1    g567(.A(G1384), .ZN(new_n993));
  AND2_X1   g568(.A1(new_n509), .A2(KEYINPUT4), .ZN(new_n994));
  INV_X1    g569(.A(new_n504), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n995), .B1(new_n481), .B2(new_n484), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n522), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n515), .A2(new_n517), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n993), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n999), .A2(new_n1000), .A3(KEYINPUT50), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT50), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT109), .B1(new_n957), .B2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(KEYINPUT108), .B(KEYINPUT50), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n957), .A2(new_n1004), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n1001), .A2(new_n1003), .A3(new_n987), .A4(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n992), .B1(new_n1006), .B2(G2084), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G8), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  NOR2_X1   g584(.A1(G168), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1008), .A2(KEYINPUT51), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1013), .B(G8), .C1(new_n1007), .C2(G286), .ZN(new_n1014));
  AOI21_X1  g589(.A(KEYINPUT120), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1007), .A2(KEYINPUT120), .A3(new_n1010), .ZN(new_n1016));
  OAI211_X1 g591(.A(new_n1012), .B(new_n1014), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  AND2_X1   g592(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1017), .A2(KEYINPUT62), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n958), .B1(new_n999), .B2(new_n988), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n990), .A2(KEYINPUT107), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT107), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n523), .A2(new_n1023), .A3(new_n989), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1021), .A2(new_n744), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G1961), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n1020), .A2(new_n1025), .B1(new_n1006), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT122), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(new_n991), .B2(G2078), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1021), .A2(KEYINPUT122), .A3(new_n744), .A4(new_n990), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(KEYINPUT53), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(G301), .B1(new_n1027), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n1009), .B1(new_n987), .B2(new_n957), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n594), .A2(G1976), .A3(new_n596), .ZN(new_n1036));
  INV_X1    g611(.A(G1976), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT52), .B1(G288), .B2(new_n1037), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1034), .A2(new_n1035), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  OAI211_X1 g614(.A(G8), .B(new_n1036), .C1(new_n999), .C2(new_n958), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1041), .B1(new_n804), .B2(G1976), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT111), .B1(new_n1040), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1040), .A2(KEYINPUT52), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n600), .A2(new_n602), .A3(G1981), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(G1981), .B1(new_n600), .B2(new_n602), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT112), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(KEYINPUT49), .ZN(new_n1049));
  INV_X1    g624(.A(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1046), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1047), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1049), .B1(new_n1052), .B2(new_n1045), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1034), .A2(new_n1051), .A3(new_n1053), .ZN(new_n1054));
  AND4_X1   g629(.A1(new_n1039), .A2(new_n1043), .A3(new_n1044), .A4(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G303), .A2(G8), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1056), .B(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n989), .ZN(new_n1060));
  AOI211_X1 g635(.A(KEYINPUT107), .B(new_n1060), .C1(new_n956), .C2(new_n518), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1023), .B1(new_n523), .B2(new_n989), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  AOI21_X1  g638(.A(G1971), .B1(new_n1063), .B2(new_n1021), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n958), .A2(G2090), .ZN(new_n1065));
  AND4_X1   g640(.A1(new_n1001), .A2(new_n1003), .A3(new_n1005), .A4(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(G8), .B(new_n1059), .C1(new_n1064), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G1971), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n987), .B1(KEYINPUT45), .B2(new_n957), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1068), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OR2_X1    g646(.A1(new_n957), .A2(new_n1004), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n523), .A2(new_n1002), .A3(new_n993), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1072), .A2(new_n776), .A3(new_n987), .A4(new_n1073), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1009), .B1(new_n1071), .B2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g650(.A(new_n1055), .B(new_n1067), .C1(new_n1059), .C2(new_n1075), .ZN(new_n1076));
  NOR4_X1   g651(.A1(new_n1018), .A2(new_n1019), .A3(new_n1033), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT124), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1007), .A2(G8), .A3(G168), .ZN(new_n1079));
  OAI21_X1  g654(.A(KEYINPUT115), .B1(new_n1076), .B2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT63), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1043), .A2(new_n1039), .A3(new_n1044), .A4(new_n1054), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1073), .B(new_n987), .C1(new_n957), .C2(new_n1004), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1083), .A2(G2090), .ZN(new_n1084));
  OAI21_X1  g659(.A(G8), .B1(new_n1064), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1082), .B1(new_n1058), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1079), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT115), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .A4(new_n1067), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1080), .A2(new_n1081), .A3(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(G8), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1059), .B1(new_n1091), .B2(KEYINPUT116), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n1092), .B1(KEYINPUT116), .B2(new_n1091), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1055), .A2(KEYINPUT113), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1082), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1067), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1098), .A2(new_n1081), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n1093), .A2(new_n1097), .A3(new_n1087), .A4(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1090), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1054), .A2(new_n1037), .A3(new_n804), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1103), .A2(new_n1046), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n1034), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1102), .A2(KEYINPUT114), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1067), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1105), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1107), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1106), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1101), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1006), .A2(new_n769), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n999), .A2(new_n958), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(new_n793), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n619), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT56), .B(G2072), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1021), .A2(new_n1022), .A3(new_n1024), .A4(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1083), .A2(new_n781), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n575), .A2(KEYINPUT57), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n582), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1123), .B1(new_n586), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(KEYINPUT117), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n1127));
  OAI211_X1 g702(.A(new_n1123), .B(new_n1127), .C1(new_n586), .C2(new_n1124), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1121), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1117), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT118), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1129), .A2(new_n1119), .A3(new_n1120), .A4(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1132), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT61), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1140), .B1(new_n1121), .B2(new_n1130), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(new_n1133), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1021), .A2(new_n961), .A3(new_n1022), .A4(new_n1024), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT119), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1063), .A2(KEYINPUT119), .A3(new_n961), .A4(new_n1021), .ZN(new_n1146));
  XOR2_X1   g721(.A(KEYINPUT58), .B(G1341), .Z(new_n1147));
  OAI21_X1  g722(.A(new_n1147), .B1(new_n999), .B2(new_n958), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1145), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(KEYINPUT59), .A3(new_n565), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1142), .A2(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1113), .A2(KEYINPUT60), .A3(new_n618), .A4(new_n1115), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1148), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1153), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n844), .B1(new_n1154), .B2(new_n1146), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1152), .B1(new_n1155), .B2(KEYINPUT59), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1151), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1116), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1113), .A2(KEYINPUT60), .A3(new_n1115), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n619), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1139), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1006), .A2(new_n1026), .ZN(new_n1163));
  NAND2_X1  g738(.A1(new_n1025), .A2(new_n1020), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1031), .A2(G301), .A3(new_n1163), .A4(new_n1164), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1165), .A2(KEYINPUT54), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1063), .A2(KEYINPUT53), .A3(new_n744), .A4(new_n1021), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1164), .A2(new_n1163), .A3(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT123), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT123), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1164), .A2(new_n1163), .A3(new_n1170), .A4(new_n1167), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1169), .A2(G171), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1166), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1134), .A2(new_n1140), .A3(new_n1136), .ZN(new_n1174));
  AND3_X1   g749(.A1(new_n1174), .A2(new_n1086), .A3(new_n1067), .ZN(new_n1175));
  XNOR2_X1  g750(.A(KEYINPUT121), .B(KEYINPUT54), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1168), .A2(G171), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1176), .B1(new_n1177), .B2(new_n1032), .ZN(new_n1178));
  NAND4_X1  g753(.A1(new_n1173), .A2(new_n1175), .A3(new_n1017), .A4(new_n1178), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1162), .A2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1078), .B1(new_n1112), .B2(new_n1180), .ZN(new_n1181));
  AOI22_X1  g756(.A1(new_n1155), .A2(KEYINPUT59), .B1(new_n1141), .B2(new_n1133), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1149), .A2(new_n565), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT59), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NAND4_X1  g760(.A1(new_n1182), .A2(new_n1161), .A3(new_n1185), .A4(new_n1152), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1186), .A2(new_n1138), .ZN(new_n1187));
  AND2_X1   g762(.A1(new_n1175), .A2(new_n1178), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1187), .A2(new_n1188), .A3(new_n1017), .A4(new_n1173), .ZN(new_n1189));
  AOI22_X1  g764(.A1(new_n1090), .A2(new_n1100), .B1(new_n1106), .B2(new_n1110), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1189), .A2(new_n1190), .A3(KEYINPUT124), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1077), .B1(new_n1181), .B2(new_n1191), .ZN(new_n1192));
  AND2_X1   g767(.A1(G290), .A2(G1986), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n959), .B1(new_n1193), .B2(new_n978), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n977), .A2(new_n1194), .ZN(new_n1195));
  XOR2_X1   g770(.A(new_n1195), .B(KEYINPUT106), .Z(new_n1196));
  OAI21_X1  g771(.A(new_n986), .B1(new_n1192), .B2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g772(.A1(G401), .A2(G227), .A3(new_n460), .ZN(new_n1199));
  NAND2_X1  g773(.A1(new_n697), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g774(.A(new_n1200), .B1(new_n946), .B2(new_n950), .ZN(new_n1201));
  AND3_X1   g775(.A1(new_n898), .A2(KEYINPUT127), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g776(.A(KEYINPUT127), .B1(new_n898), .B2(new_n1201), .ZN(new_n1203));
  NOR2_X1   g777(.A1(new_n1202), .A2(new_n1203), .ZN(G308));
  NAND2_X1  g778(.A1(new_n898), .A2(new_n1201), .ZN(new_n1205));
  INV_X1    g779(.A(KEYINPUT127), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g781(.A1(new_n898), .A2(KEYINPUT127), .A3(new_n1201), .ZN(new_n1208));
  NAND2_X1  g782(.A1(new_n1207), .A2(new_n1208), .ZN(G225));
endmodule


