//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n973,
    new_n974, new_n975, new_n976, new_n978, new_n979, new_n980, new_n981,
    new_n982;
  XNOR2_X1  g000(.A(G197gat), .B(G204gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT22), .ZN(new_n203));
  INV_X1    g002(.A(G211gat), .ZN(new_n204));
  INV_X1    g003(.A(G218gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n208), .A2(new_n202), .A3(new_n206), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n210), .A2(KEYINPUT70), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT70), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n207), .A2(new_n213), .A3(new_n209), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G183gat), .ZN(new_n216));
  INV_X1    g015(.A(G190gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT24), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT64), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n221), .A2(new_n224), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n218), .B(new_n223), .C1(new_n225), .C2(new_n222), .ZN(new_n226));
  NAND2_X1  g025(.A1(G169gat), .A2(G176gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT23), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n226), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT25), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n227), .B(KEYINPUT65), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n221), .A2(new_n218), .A3(new_n224), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n230), .A2(KEYINPUT25), .A3(new_n234), .A4(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n236), .A2(new_n237), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n233), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(G226gat), .ZN(new_n241));
  INV_X1    g040(.A(G233gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT28), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT27), .B(G183gat), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(KEYINPUT67), .ZN(new_n247));
  AND2_X1   g046(.A1(new_n216), .A2(KEYINPUT27), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT67), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n217), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n245), .B1(new_n247), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n246), .A2(KEYINPUT28), .A3(new_n217), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n251), .A2(new_n252), .B1(G183gat), .B2(G190gat), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT26), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n228), .A2(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n227), .A3(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  AND3_X1   g057(.A1(new_n240), .A2(new_n244), .A3(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n243), .A2(KEYINPUT29), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n260), .B1(new_n240), .B2(new_n258), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n215), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n240), .A2(new_n244), .A3(new_n258), .ZN(new_n263));
  INV_X1    g062(.A(new_n215), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n236), .B(KEYINPUT66), .ZN(new_n265));
  AOI22_X1  g064(.A1(new_n265), .A2(new_n233), .B1(new_n253), .B2(new_n257), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n263), .B(new_n264), .C1(new_n260), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT30), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n262), .A2(KEYINPUT30), .A3(new_n267), .ZN(new_n271));
  XNOR2_X1  g070(.A(G8gat), .B(G36gat), .ZN(new_n272));
  INV_X1    g071(.A(G64gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n272), .B(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G92gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n270), .A2(new_n271), .A3(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(G120gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G113gat), .ZN(new_n280));
  INV_X1    g079(.A(G113gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G120gat), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT1), .B1(new_n280), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G127gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G134gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G141gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(G148gat), .ZN(new_n289));
  XNOR2_X1  g088(.A(KEYINPUT71), .B(G148gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n289), .B1(new_n290), .B2(new_n288), .ZN(new_n291));
  NAND2_X1  g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292));
  INV_X1    g091(.A(G155gat), .ZN(new_n293));
  INV_X1    g092(.A(G162gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n292), .B1(new_n295), .B2(KEYINPUT2), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n291), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G141gat), .B(G148gat), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n292), .B(new_n295), .C1(new_n298), .C2(KEYINPUT2), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  OR2_X1    g099(.A1(new_n283), .A2(new_n284), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n283), .A2(new_n284), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(G134gat), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT4), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT4), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n287), .A2(new_n300), .A3(new_n306), .A4(new_n303), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n287), .A2(new_n303), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n297), .A2(new_n299), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT3), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT73), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT72), .B(KEYINPUT3), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n312), .B1(new_n300), .B2(new_n313), .ZN(new_n314));
  NAND4_X1  g113(.A1(new_n297), .A2(new_n312), .A3(new_n299), .A4(new_n313), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n309), .B(new_n311), .C1(new_n314), .C2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G225gat), .A2(G233gat), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n308), .A2(new_n317), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT5), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n309), .A2(new_n310), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(new_n304), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n322), .B1(new_n324), .B2(new_n319), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n313), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT73), .B1(new_n310), .B2(new_n327), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n328), .A2(new_n315), .B1(new_n303), .B2(new_n287), .ZN(new_n329));
  AOI22_X1  g128(.A1(new_n311), .A2(new_n329), .B1(new_n305), .B2(new_n307), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n319), .A2(KEYINPUT5), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(G1gat), .B(G29gat), .Z(new_n334));
  XNOR2_X1  g133(.A(G57gat), .B(G85gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT74), .B(KEYINPUT0), .ZN(new_n337));
  XOR2_X1   g136(.A(new_n336), .B(new_n337), .Z(new_n338));
  NAND2_X1  g137(.A1(new_n333), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g138(.A1(new_n262), .A2(KEYINPUT30), .A3(new_n267), .A4(new_n276), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n318), .B1(new_n308), .B2(new_n317), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT39), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n338), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n323), .A2(new_n318), .A3(new_n304), .ZN(new_n344));
  OAI211_X1 g143(.A(KEYINPUT39), .B(new_n344), .C1(new_n330), .C2(new_n318), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(new_n345), .A3(KEYINPUT40), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n278), .A2(new_n339), .A3(new_n340), .A4(new_n346), .ZN(new_n347));
  AOI21_X1  g146(.A(KEYINPUT40), .B1(new_n343), .B2(new_n345), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n215), .A2(KEYINPUT29), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n310), .B1(new_n350), .B2(KEYINPUT3), .ZN(new_n351));
  AND2_X1   g150(.A1(G228gat), .A2(G233gat), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT29), .B1(new_n328), .B2(new_n315), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n351), .B(new_n352), .C1(new_n264), .C2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n210), .A2(KEYINPUT75), .A3(new_n211), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT29), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n355), .B(new_n356), .C1(KEYINPUT75), .C2(new_n211), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n300), .B1(new_n357), .B2(new_n313), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n356), .B1(new_n314), .B2(new_n316), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(new_n215), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n354), .B1(new_n360), .B2(new_n352), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(G22gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT31), .ZN(new_n364));
  INV_X1    g163(.A(G50gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT76), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n362), .A2(new_n368), .ZN(new_n369));
  OR2_X1    g168(.A1(new_n361), .A2(G22gat), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n361), .A2(G22gat), .A3(new_n367), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n369), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT77), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n361), .A2(G22gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n374), .A2(new_n366), .ZN(new_n375));
  AND3_X1   g174(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n373), .B1(new_n372), .B2(new_n375), .ZN(new_n377));
  NOR3_X1   g176(.A1(new_n349), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT6), .ZN(new_n379));
  AOI22_X1  g178(.A1(new_n321), .A2(new_n325), .B1(new_n330), .B2(new_n331), .ZN(new_n380));
  INV_X1    g179(.A(new_n338), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n339), .A2(new_n379), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT79), .B(KEYINPUT38), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT37), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n262), .A2(new_n385), .A3(new_n267), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n385), .B1(new_n262), .B2(new_n267), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n384), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT80), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n381), .B1(new_n326), .B2(new_n332), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n390), .B1(new_n391), .B2(KEYINPUT6), .ZN(new_n392));
  NOR4_X1   g191(.A1(new_n380), .A2(KEYINPUT80), .A3(new_n379), .A4(new_n381), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n383), .B(new_n389), .C1(new_n392), .C2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n384), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n268), .A2(new_n277), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT78), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n262), .A2(new_n398), .A3(new_n267), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n259), .A2(new_n261), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(KEYINPUT78), .A3(new_n264), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(KEYINPUT37), .A3(new_n401), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n402), .A2(new_n396), .A3(new_n386), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n397), .B1(new_n403), .B2(new_n277), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n395), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT36), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT68), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n240), .A2(new_n258), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n309), .ZN(new_n409));
  INV_X1    g208(.A(new_n309), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n266), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(G227gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(new_n242), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n407), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n414), .ZN(new_n416));
  AOI211_X1 g215(.A(KEYINPUT68), .B(new_n416), .C1(new_n409), .C2(new_n411), .ZN(new_n417));
  OAI21_X1  g216(.A(KEYINPUT32), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n409), .A2(new_n416), .A3(new_n411), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT34), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT34), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n409), .A2(new_n411), .A3(new_n421), .A4(new_n416), .ZN(new_n422));
  AND2_X1   g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT69), .B(G71gat), .ZN(new_n425));
  INV_X1    g224(.A(G99gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(new_n425), .B(new_n426), .ZN(new_n427));
  XNOR2_X1  g226(.A(G15gat), .B(G43gat), .ZN(new_n428));
  XOR2_X1   g227(.A(new_n427), .B(new_n428), .Z(new_n429));
  INV_X1    g228(.A(new_n429), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n240), .A2(new_n410), .A3(new_n258), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n410), .B1(new_n240), .B2(new_n258), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n414), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT68), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n412), .A2(new_n407), .A3(new_n414), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT33), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n430), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n420), .A2(new_n422), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n436), .A2(new_n439), .A3(KEYINPUT32), .ZN(new_n440));
  AND3_X1   g239(.A1(new_n424), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n438), .B1(new_n424), .B2(new_n440), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n406), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n436), .A2(new_n437), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(new_n429), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n418), .A2(new_n423), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n439), .B1(new_n436), .B2(KEYINPUT32), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n424), .A2(new_n438), .A3(new_n440), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(KEYINPUT36), .A3(new_n449), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n378), .A2(new_n405), .B1(new_n443), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n391), .A2(KEYINPUT6), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n383), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n278), .A2(new_n340), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n455), .B1(new_n376), .B2(new_n377), .ZN(new_n456));
  AND3_X1   g255(.A1(new_n361), .A2(G22gat), .A3(new_n367), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n367), .B1(new_n361), .B2(G22gat), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n457), .A2(new_n458), .A3(new_n374), .ZN(new_n459));
  INV_X1    g258(.A(new_n375), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT77), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n372), .A2(new_n373), .A3(new_n375), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n461), .A2(new_n448), .A3(new_n462), .A4(new_n449), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT35), .B1(new_n463), .B2(new_n455), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n376), .A2(new_n377), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n441), .A2(new_n442), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n383), .B1(new_n392), .B2(new_n393), .ZN(new_n467));
  XOR2_X1   g266(.A(KEYINPUT81), .B(KEYINPUT35), .Z(new_n468));
  AND3_X1   g267(.A1(new_n467), .A2(new_n454), .A3(new_n468), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n465), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n451), .A2(new_n456), .B1(new_n464), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G29gat), .A2(G36gat), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  OR2_X1    g272(.A1(KEYINPUT84), .A2(G43gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(KEYINPUT84), .A2(G43gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n474), .A2(new_n365), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n365), .A2(G43gat), .ZN(new_n477));
  INV_X1    g276(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT15), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n473), .B1(new_n479), .B2(KEYINPUT85), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT85), .ZN(new_n481));
  AND2_X1   g280(.A1(KEYINPUT84), .A2(G43gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(KEYINPUT84), .A2(G43gat), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n477), .B1(new_n484), .B2(new_n365), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n481), .B1(new_n485), .B2(KEYINPUT15), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n365), .A2(G43gat), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n478), .A2(KEYINPUT15), .A3(new_n487), .ZN(new_n488));
  NOR3_X1   g287(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n480), .A2(new_n486), .A3(new_n488), .A4(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT82), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT83), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n491), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n495), .B1(new_n491), .B2(new_n494), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n490), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n491), .A2(new_n494), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(KEYINPUT83), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n491), .A2(new_n494), .A3(new_n495), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n489), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n498), .A2(new_n502), .A3(new_n472), .ZN(new_n503));
  INV_X1    g302(.A(new_n488), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n493), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(G15gat), .B(G22gat), .Z(new_n507));
  INV_X1    g306(.A(G1gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(G15gat), .B(G22gat), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT16), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(G1gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT86), .ZN(new_n514));
  INV_X1    g313(.A(G8gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n515), .ZN(new_n517));
  NAND2_X1  g316(.A1(KEYINPUT86), .A2(G8gat), .ZN(new_n518));
  NAND4_X1  g317(.A1(new_n509), .A2(new_n512), .A3(new_n517), .A4(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n506), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(G229gat), .A2(G233gat), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n493), .A2(new_n505), .A3(KEYINPUT17), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n516), .A2(new_n519), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT17), .B1(new_n493), .B2(new_n505), .ZN(new_n525));
  OAI211_X1 g324(.A(new_n520), .B(new_n521), .C1(new_n524), .C2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(KEYINPUT87), .A2(KEYINPUT18), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g327(.A(new_n521), .B(KEYINPUT13), .Z(new_n529));
  INV_X1    g328(.A(new_n520), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n506), .B1(new_n516), .B2(new_n519), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT17), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n506), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(new_n523), .A3(new_n522), .ZN(new_n535));
  INV_X1    g334(.A(new_n527), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n535), .A2(new_n520), .A3(new_n521), .A4(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n528), .A2(new_n532), .A3(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT11), .B(G169gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(G197gat), .ZN(new_n540));
  XOR2_X1   g339(.A(G113gat), .B(G141gat), .Z(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT12), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n538), .A2(new_n544), .ZN(new_n545));
  NAND4_X1  g344(.A1(new_n528), .A2(new_n537), .A3(new_n543), .A4(new_n532), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT88), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n471), .A2(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n551));
  XNOR2_X1  g350(.A(G183gat), .B(G211gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT21), .ZN(new_n555));
  AND2_X1   g354(.A1(G71gat), .A2(G78gat), .ZN(new_n556));
  NOR2_X1   g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  XNOR2_X1  g357(.A(G57gat), .B(G64gat), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT9), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G71gat), .ZN(new_n562));
  INV_X1    g361(.A(G78gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g363(.A1(G71gat), .A2(G78gat), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT89), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n273), .A2(G57gat), .ZN(new_n568));
  INV_X1    g367(.A(G57gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(G64gat), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  AND3_X1   g370(.A1(new_n566), .A2(new_n567), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n567), .B1(new_n566), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n561), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n523), .B1(new_n555), .B2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n575), .B(KEYINPUT91), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT90), .B(KEYINPUT21), .Z(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n578), .B(KEYINPUT92), .ZN(new_n579));
  OR2_X1    g378(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n579), .ZN(new_n581));
  XNOR2_X1  g380(.A(G127gat), .B(G155gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n582), .B(new_n583), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n580), .A2(new_n581), .A3(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n585), .B1(new_n580), .B2(new_n581), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n554), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n590), .A2(new_n553), .A3(new_n586), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G190gat), .B(G218gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(new_n286), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT95), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(KEYINPUT95), .A2(G99gat), .A3(G106gat), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n597), .A2(KEYINPUT8), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n275), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n600));
  OAI21_X1  g399(.A(G92gat), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n601));
  AND2_X1   g400(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G99gat), .B(G106gat), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n599), .A2(new_n603), .A3(new_n605), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n534), .A2(new_n609), .A3(new_n522), .ZN(new_n610));
  NAND3_X1  g409(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n611));
  INV_X1    g410(.A(new_n506), .ZN(new_n612));
  OAI211_X1 g411(.A(new_n610), .B(new_n611), .C1(new_n612), .C2(new_n609), .ZN(new_n613));
  AOI21_X1  g412(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n594), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n613), .A2(new_n614), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n613), .A2(new_n614), .ZN(new_n619));
  INV_X1    g418(.A(new_n594), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g421(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(G162gat), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n617), .A2(new_n621), .A3(new_n624), .ZN(new_n627));
  XNOR2_X1  g426(.A(G176gat), .B(G204gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT97), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(G120gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G148gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(G230gat), .A2(G233gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n632), .B(KEYINPUT98), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n609), .A2(new_n574), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n556), .B1(KEYINPUT9), .B2(new_n557), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT89), .B1(new_n637), .B2(new_n559), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n566), .A2(new_n567), .A3(new_n571), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n640), .A2(new_n561), .A3(new_n608), .A4(new_n607), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n635), .A2(new_n636), .A3(new_n641), .ZN(new_n642));
  AND2_X1   g441(.A1(new_n607), .A2(new_n608), .ZN(new_n643));
  NAND4_X1  g442(.A1(new_n643), .A2(KEYINPUT10), .A3(new_n640), .A4(new_n561), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n634), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n632), .B1(new_n635), .B2(new_n641), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n631), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(KEYINPUT99), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(KEYINPUT96), .ZN(new_n649));
  INV_X1    g448(.A(G148gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n630), .B(new_n650), .ZN(new_n651));
  AOI22_X1  g450(.A1(new_n642), .A2(new_n644), .B1(G230gat), .B2(G233gat), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT96), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(new_n649), .B(new_n651), .C1(new_n654), .C2(new_n646), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n648), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND4_X1  g456(.A1(new_n592), .A2(new_n626), .A3(new_n627), .A4(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n550), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n660), .A2(new_n453), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(new_n508), .ZN(G1324gat));
  NOR2_X1   g461(.A1(new_n660), .A2(new_n454), .ZN(new_n663));
  NAND2_X1  g462(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n511), .A2(new_n515), .ZN(new_n665));
  AND3_X1   g464(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n666), .A2(KEYINPUT42), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(KEYINPUT42), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n667), .B(new_n668), .C1(new_n515), .C2(new_n663), .ZN(G1325gat));
  INV_X1    g468(.A(G15gat), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n443), .A2(new_n450), .ZN(new_n671));
  NOR3_X1   g470(.A1(new_n660), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n550), .A2(new_n659), .A3(new_n466), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n672), .B1(new_n670), .B2(new_n673), .ZN(G1326gat));
  NOR2_X1   g473(.A1(new_n660), .A2(new_n465), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT43), .B(G22gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  AND2_X1   g476(.A1(new_n626), .A2(new_n627), .ZN(new_n678));
  NOR3_X1   g477(.A1(new_n678), .A2(new_n592), .A3(new_n656), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n550), .A2(new_n679), .ZN(new_n680));
  NOR3_X1   g479(.A1(new_n680), .A2(G29gat), .A3(new_n453), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT45), .Z(new_n682));
  OAI21_X1  g481(.A(KEYINPUT44), .B1(new_n471), .B2(new_n678), .ZN(new_n683));
  INV_X1    g482(.A(new_n349), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n405), .A2(new_n465), .A3(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n456), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g486(.A(KEYINPUT101), .B(new_n455), .C1(new_n376), .C2(new_n377), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n685), .A2(new_n687), .A3(new_n671), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n464), .A2(new_n470), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n626), .A2(new_n627), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT102), .B(KEYINPUT44), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n656), .B1(new_n683), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT100), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n592), .B(new_n697), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n698), .A2(new_n547), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n453), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n682), .A2(new_n701), .ZN(G1328gat));
  AND2_X1   g501(.A1(new_n550), .A2(new_n679), .ZN(new_n703));
  INV_X1    g502(.A(G36gat), .ZN(new_n704));
  INV_X1    g503(.A(new_n454), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n706), .A2(KEYINPUT46), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT103), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n706), .A2(KEYINPUT46), .ZN(new_n710));
  OAI21_X1  g509(.A(G36gat), .B1(new_n700), .B2(new_n454), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n709), .A2(new_n710), .A3(new_n711), .ZN(G1329gat));
  OAI21_X1  g511(.A(new_n484), .B1(new_n700), .B2(new_n671), .ZN(new_n713));
  INV_X1    g512(.A(new_n466), .ZN(new_n714));
  OR3_X1    g513(.A1(new_n680), .A2(new_n484), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT47), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1330gat));
  OAI21_X1  g517(.A(KEYINPUT104), .B1(new_n700), .B2(new_n465), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT104), .ZN(new_n720));
  INV_X1    g519(.A(new_n465), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n696), .A2(new_n720), .A3(new_n721), .A4(new_n699), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n719), .A2(G50gat), .A3(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n703), .A2(new_n365), .A3(new_n721), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n723), .A2(KEYINPUT48), .A3(new_n724), .ZN(new_n725));
  OAI21_X1  g524(.A(G50gat), .B1(new_n700), .B2(new_n465), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n724), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT48), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n725), .A2(new_n729), .ZN(G1331gat));
  AOI21_X1  g529(.A(new_n547), .B1(new_n689), .B2(new_n690), .ZN(new_n731));
  INV_X1    g530(.A(new_n592), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n692), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n731), .A2(new_n733), .A3(new_n656), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n453), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(new_n569), .ZN(G1332gat));
  INV_X1    g535(.A(new_n734), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n454), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT105), .Z(new_n740));
  NOR2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(G1333gat));
  OAI21_X1  g541(.A(new_n562), .B1(new_n734), .B2(new_n714), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n737), .A2(G71gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(new_n671), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g545(.A1(new_n734), .A2(new_n465), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(new_n563), .ZN(G1335gat));
  NOR2_X1   g547(.A1(new_n657), .A2(new_n547), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  AOI211_X1 g549(.A(new_n592), .B(new_n750), .C1(new_n683), .C2(new_n695), .ZN(new_n751));
  INV_X1    g550(.A(new_n453), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n751), .A2(G85gat), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT51), .ZN(new_n754));
  INV_X1    g553(.A(new_n547), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n678), .A2(new_n592), .ZN(new_n756));
  AND4_X1   g555(.A1(new_n754), .A2(new_n691), .A3(new_n755), .A4(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n754), .B1(new_n731), .B2(new_n756), .ZN(new_n758));
  NOR4_X1   g557(.A1(new_n757), .A2(new_n758), .A3(new_n453), .A4(new_n657), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n753), .B1(G85gat), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n760), .B(new_n761), .ZN(G1336gat));
  INV_X1    g561(.A(KEYINPUT52), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n275), .B1(new_n751), .B2(new_n705), .ZN(new_n764));
  INV_X1    g563(.A(KEYINPUT107), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n763), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NOR2_X1   g565(.A1(new_n757), .A2(new_n758), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n767), .A2(new_n275), .A3(new_n656), .A4(new_n705), .ZN(new_n768));
  AOI211_X1 g567(.A(new_n678), .B(new_n693), .C1(new_n689), .C2(new_n690), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT44), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n685), .A2(new_n671), .A3(new_n456), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n690), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n770), .B1(new_n772), .B2(new_n692), .ZN(new_n773));
  OAI211_X1 g572(.A(new_n732), .B(new_n749), .C1(new_n769), .C2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G92gat), .B1(new_n774), .B2(new_n454), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT108), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n768), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n776), .B1(new_n768), .B2(new_n775), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n766), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n691), .A2(new_n755), .A3(new_n756), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT51), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n731), .A2(new_n754), .A3(new_n756), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n781), .A2(new_n275), .A3(new_n656), .A4(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(new_n454), .ZN(new_n784));
  OAI21_X1  g583(.A(KEYINPUT108), .B1(new_n764), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(KEYINPUT52), .B1(new_n775), .B2(KEYINPUT107), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n768), .A2(new_n775), .A3(new_n776), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n779), .A2(new_n788), .ZN(G1337gat));
  OAI21_X1  g588(.A(G99gat), .B1(new_n774), .B2(new_n671), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n767), .A2(new_n426), .A3(new_n656), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n791), .B2(new_n714), .ZN(G1338gat));
  INV_X1    g591(.A(G106gat), .ZN(new_n793));
  AND4_X1   g592(.A1(new_n793), .A2(new_n767), .A3(new_n656), .A4(new_n721), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n751), .B2(new_n721), .ZN(new_n795));
  OR3_X1    g594(.A1(new_n794), .A2(new_n795), .A3(KEYINPUT53), .ZN(new_n796));
  OAI21_X1  g595(.A(KEYINPUT53), .B1(new_n794), .B2(new_n795), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(G1339gat));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n800), .B1(new_n659), .B2(new_n755), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n658), .A2(KEYINPUT109), .A3(new_n547), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n530), .A2(new_n531), .A3(new_n529), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n521), .B1(new_n535), .B2(new_n520), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n542), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n546), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n656), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n642), .A2(new_n644), .A3(new_n634), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n652), .ZN(new_n810));
  AOI211_X1 g609(.A(KEYINPUT54), .B(new_n634), .C1(new_n642), .C2(new_n644), .ZN(new_n811));
  OAI21_X1  g610(.A(KEYINPUT110), .B1(new_n811), .B2(new_n651), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n642), .A2(new_n644), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n813), .A2(new_n814), .A3(new_n633), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT110), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n816), .A3(new_n631), .ZN(new_n817));
  AOI221_X4 g616(.A(KEYINPUT55), .B1(new_n810), .B2(KEYINPUT54), .C1(new_n812), .C2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT55), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n812), .A2(new_n817), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n810), .A2(KEYINPUT54), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n655), .B1(new_n818), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n808), .B1(new_n823), .B2(new_n755), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT111), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n547), .B(new_n655), .C1(new_n822), .C2(new_n818), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT111), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n827), .A3(new_n808), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n825), .A2(new_n678), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT112), .ZN(new_n830));
  INV_X1    g629(.A(new_n823), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n692), .A2(new_n831), .A3(new_n807), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n698), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n830), .B1(new_n829), .B2(new_n832), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n803), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n463), .A2(new_n453), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n836), .A2(KEYINPUT114), .A3(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT114), .B1(new_n836), .B2(new_n837), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n839), .A2(new_n840), .A3(new_n705), .ZN(new_n841));
  AOI21_X1  g640(.A(G113gat), .B1(new_n841), .B2(new_n547), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n705), .A2(new_n453), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT113), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n826), .A2(new_n827), .A3(new_n808), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n827), .B1(new_n826), .B2(new_n808), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n845), .A2(new_n846), .A3(new_n692), .ZN(new_n847));
  INV_X1    g646(.A(new_n832), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT112), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n849), .A2(new_n698), .A3(new_n833), .ZN(new_n850));
  AOI211_X1 g649(.A(new_n844), .B(new_n721), .C1(new_n850), .C2(new_n803), .ZN(new_n851));
  AOI21_X1  g650(.A(KEYINPUT113), .B1(new_n836), .B2(new_n465), .ZN(new_n852));
  OAI211_X1 g651(.A(new_n466), .B(new_n843), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(new_n281), .A3(new_n549), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n799), .B1(new_n842), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n840), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n856), .A2(new_n454), .A3(new_n838), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n281), .B1(new_n857), .B2(new_n755), .ZN(new_n858));
  INV_X1    g657(.A(new_n852), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n721), .B1(new_n850), .B2(new_n803), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n860), .A2(KEYINPUT113), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n862), .A2(G113gat), .A3(new_n466), .A4(new_n843), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n858), .B(KEYINPUT115), .C1(new_n863), .C2(new_n549), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n855), .A2(new_n864), .ZN(G1340gat));
  NAND3_X1  g664(.A1(new_n841), .A2(new_n279), .A3(new_n656), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n862), .A2(new_n656), .A3(new_n466), .A4(new_n843), .ZN(new_n867));
  AOI21_X1  g666(.A(KEYINPUT116), .B1(new_n867), .B2(G120gat), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT116), .B(G120gat), .C1(new_n853), .C2(new_n657), .ZN(new_n869));
  INV_X1    g668(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n866), .B1(new_n868), .B2(new_n870), .ZN(G1341gat));
  AOI21_X1  g670(.A(G127gat), .B1(new_n841), .B2(new_n592), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n853), .A2(new_n284), .A3(new_n698), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n872), .A2(new_n873), .ZN(G1342gat));
  NOR2_X1   g673(.A1(new_n678), .A2(G134gat), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n856), .A2(new_n454), .A3(new_n838), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(KEYINPUT117), .ZN(new_n878));
  OR2_X1    g677(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n879));
  OAI21_X1  g678(.A(G134gat), .B1(new_n853), .B2(new_n678), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n876), .A2(new_n881), .A3(KEYINPUT56), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n878), .A2(new_n879), .A3(new_n880), .A4(new_n882), .ZN(G1343gat));
  AND2_X1   g682(.A1(new_n671), .A2(new_n843), .ZN(new_n884));
  XOR2_X1   g683(.A(new_n884), .B(KEYINPUT118), .Z(new_n885));
  AOI21_X1  g684(.A(new_n465), .B1(new_n850), .B2(new_n803), .ZN(new_n886));
  XOR2_X1   g685(.A(KEYINPUT119), .B(KEYINPUT57), .Z(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT57), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n548), .A2(new_n831), .B1(new_n656), .B2(new_n807), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n832), .B1(new_n890), .B2(new_n692), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n732), .ZN(new_n892));
  AOI211_X1 g691(.A(new_n889), .B(new_n465), .C1(new_n803), .C2(new_n892), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n885), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n288), .B1(new_n895), .B2(new_n548), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n886), .A2(new_n884), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n548), .A2(KEYINPUT120), .A3(new_n288), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT120), .B1(new_n548), .B2(new_n288), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n900), .A2(KEYINPUT58), .ZN(new_n901));
  OAI211_X1 g700(.A(new_n547), .B(new_n885), .C1(new_n888), .C2(new_n893), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n900), .B1(new_n902), .B2(G141gat), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT58), .ZN(new_n904));
  OAI22_X1  g703(.A1(new_n896), .A2(new_n901), .B1(new_n903), .B2(new_n904), .ZN(G1344gat));
  NOR3_X1   g704(.A1(new_n897), .A2(new_n290), .A3(new_n657), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT121), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n656), .B(new_n885), .C1(new_n888), .C2(new_n893), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT59), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n908), .A2(new_n909), .A3(new_n290), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n886), .A2(new_n887), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT122), .B1(new_n658), .B2(new_n548), .ZN(new_n912));
  OR3_X1    g711(.A1(new_n658), .A2(KEYINPUT122), .A3(new_n548), .ZN(new_n913));
  AND3_X1   g712(.A1(new_n892), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n889), .B1(new_n914), .B2(new_n465), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n656), .A3(new_n885), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n909), .B1(new_n917), .B2(G148gat), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n907), .B1(new_n910), .B2(new_n918), .ZN(G1345gat));
  INV_X1    g718(.A(new_n897), .ZN(new_n920));
  AOI21_X1  g719(.A(G155gat), .B1(new_n920), .B2(new_n592), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n698), .A2(new_n293), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n921), .B1(new_n895), .B2(new_n922), .ZN(G1346gat));
  AOI21_X1  g722(.A(G162gat), .B1(new_n920), .B2(new_n692), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n678), .A2(new_n294), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n895), .B2(new_n925), .ZN(G1347gat));
  NOR2_X1   g725(.A1(new_n752), .A2(new_n454), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT123), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n466), .B(new_n929), .C1(new_n851), .C2(new_n852), .ZN(new_n930));
  OAI21_X1  g729(.A(G169gat), .B1(new_n930), .B2(new_n549), .ZN(new_n931));
  AND3_X1   g730(.A1(new_n860), .A2(new_n466), .A3(new_n927), .ZN(new_n932));
  INV_X1    g731(.A(G169gat), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(new_n933), .A3(new_n547), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n931), .A2(new_n934), .ZN(G1348gat));
  AOI21_X1  g734(.A(G176gat), .B1(new_n932), .B2(new_n656), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n930), .A2(new_n657), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(G176gat), .ZN(G1349gat));
  OAI21_X1  g737(.A(G183gat), .B1(new_n930), .B2(new_n698), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n932), .A2(new_n592), .A3(new_n246), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT60), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT60), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n939), .A2(new_n943), .A3(new_n940), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n942), .A2(new_n944), .ZN(G1350gat));
  NAND3_X1  g744(.A1(new_n932), .A2(new_n217), .A3(new_n692), .ZN(new_n946));
  XNOR2_X1  g745(.A(new_n946), .B(KEYINPUT124), .ZN(new_n947));
  OAI211_X1 g746(.A(KEYINPUT61), .B(G190gat), .C1(new_n930), .C2(new_n678), .ZN(new_n948));
  OAI21_X1  g747(.A(G190gat), .B1(new_n930), .B2(new_n678), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT61), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n947), .A2(new_n948), .A3(new_n951), .ZN(G1351gat));
  AND2_X1   g751(.A1(new_n886), .A2(new_n671), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n927), .ZN(new_n954));
  INV_X1    g753(.A(new_n954), .ZN(new_n955));
  INV_X1    g754(.A(G197gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n955), .A2(new_n956), .A3(new_n547), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n929), .A2(new_n671), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT125), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n959), .B1(new_n911), .B2(new_n915), .ZN(new_n960));
  AND2_X1   g759(.A1(new_n960), .A2(new_n548), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n957), .B1(new_n961), .B2(new_n956), .ZN(G1352gat));
  INV_X1    g761(.A(new_n959), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n916), .A2(new_n656), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n964), .A2(KEYINPUT126), .ZN(new_n965));
  INV_X1    g764(.A(KEYINPUT126), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n916), .A2(new_n966), .A3(new_n656), .A4(new_n963), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n965), .A2(new_n967), .A3(G204gat), .ZN(new_n968));
  OR2_X1    g767(.A1(new_n657), .A2(G204gat), .ZN(new_n969));
  OAI21_X1  g768(.A(KEYINPUT62), .B1(new_n954), .B2(new_n969), .ZN(new_n970));
  OR3_X1    g769(.A1(new_n954), .A2(KEYINPUT62), .A3(new_n969), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(G1353gat));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n204), .A3(new_n592), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n960), .A2(new_n592), .ZN(new_n974));
  AND3_X1   g773(.A1(new_n974), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n975));
  AOI21_X1  g774(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n973), .B1(new_n975), .B2(new_n976), .ZN(G1354gat));
  NAND2_X1  g776(.A1(new_n960), .A2(KEYINPUT127), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(new_n692), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n960), .A2(KEYINPUT127), .ZN(new_n980));
  OAI21_X1  g779(.A(G218gat), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND3_X1  g780(.A1(new_n955), .A2(new_n205), .A3(new_n692), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(G1355gat));
endmodule


