

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U550 ( .A(n634), .B(n613), .ZN(n623) );
  AND2_X2 U551 ( .A1(n519), .A2(G2104), .ZN(n883) );
  NOR2_X2 U552 ( .A1(n523), .A2(n522), .ZN(G160) );
  NOR2_X1 U553 ( .A1(n632), .A2(n631), .ZN(n633) );
  INV_X1 U554 ( .A(KEYINPUT26), .ZN(n608) );
  AND2_X1 U555 ( .A1(n623), .A2(G2072), .ZN(n622) );
  INV_X1 U556 ( .A(KEYINPUT91), .ZN(n613) );
  NOR2_X1 U557 ( .A1(n675), .A2(n689), .ZN(n676) );
  XNOR2_X1 U558 ( .A(n661), .B(KEYINPUT32), .ZN(n671) );
  NOR2_X1 U559 ( .A1(n684), .A2(n683), .ZN(n691) );
  NOR2_X1 U560 ( .A1(G651), .A2(n542), .ZN(n788) );
  AND2_X1 U561 ( .A1(G2104), .A2(G2105), .ZN(n879) );
  NAND2_X1 U562 ( .A1(G113), .A2(n879), .ZN(n514) );
  XNOR2_X1 U563 ( .A(n514), .B(KEYINPUT64), .ZN(n517) );
  INV_X1 U564 ( .A(G2105), .ZN(n519) );
  NAND2_X1 U565 ( .A1(G101), .A2(n883), .ZN(n515) );
  XOR2_X1 U566 ( .A(KEYINPUT23), .B(n515), .Z(n516) );
  NAND2_X1 U567 ( .A1(n517), .A2(n516), .ZN(n523) );
  NOR2_X1 U568 ( .A1(G2104), .A2(G2105), .ZN(n518) );
  XOR2_X2 U569 ( .A(KEYINPUT17), .B(n518), .Z(n885) );
  NAND2_X1 U570 ( .A1(G137), .A2(n885), .ZN(n521) );
  NOR2_X2 U571 ( .A1(G2104), .A2(n519), .ZN(n880) );
  NAND2_X1 U572 ( .A1(G125), .A2(n880), .ZN(n520) );
  NAND2_X1 U573 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U574 ( .A1(G651), .A2(G543), .ZN(n783) );
  NAND2_X1 U575 ( .A1(G86), .A2(n783), .ZN(n528) );
  INV_X1 U576 ( .A(KEYINPUT1), .ZN(n526) );
  INV_X1 U577 ( .A(G651), .ZN(n529) );
  NOR2_X1 U578 ( .A1(G543), .A2(n529), .ZN(n524) );
  XNOR2_X1 U579 ( .A(KEYINPUT66), .B(n524), .ZN(n525) );
  XNOR2_X2 U580 ( .A(n526), .B(n525), .ZN(n789) );
  NAND2_X1 U581 ( .A1(G61), .A2(n789), .ZN(n527) );
  NAND2_X1 U582 ( .A1(n528), .A2(n527), .ZN(n532) );
  XOR2_X1 U583 ( .A(KEYINPUT0), .B(G543), .Z(n542) );
  NOR2_X1 U584 ( .A1(n542), .A2(n529), .ZN(n784) );
  NAND2_X1 U585 ( .A1(n784), .A2(G73), .ZN(n530) );
  XOR2_X1 U586 ( .A(KEYINPUT2), .B(n530), .Z(n531) );
  NOR2_X1 U587 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U588 ( .A(n533), .B(KEYINPUT80), .ZN(n535) );
  NAND2_X1 U589 ( .A1(G48), .A2(n788), .ZN(n534) );
  NAND2_X1 U590 ( .A1(n535), .A2(n534), .ZN(G305) );
  AND2_X1 U591 ( .A1(G138), .A2(n885), .ZN(n541) );
  NAND2_X1 U592 ( .A1(G102), .A2(n883), .ZN(n539) );
  NAND2_X1 U593 ( .A1(G126), .A2(n880), .ZN(n537) );
  NAND2_X1 U594 ( .A1(G114), .A2(n879), .ZN(n536) );
  AND2_X1 U595 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U596 ( .A1(n539), .A2(n538), .ZN(n540) );
  NOR2_X1 U597 ( .A1(n541), .A2(n540), .ZN(G164) );
  NAND2_X1 U598 ( .A1(G87), .A2(n542), .ZN(n544) );
  NAND2_X1 U599 ( .A1(G74), .A2(G651), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U601 ( .A1(n789), .A2(n545), .ZN(n547) );
  NAND2_X1 U602 ( .A1(n788), .A2(G49), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n547), .A2(n546), .ZN(G288) );
  NAND2_X1 U604 ( .A1(G91), .A2(n783), .ZN(n549) );
  NAND2_X1 U605 ( .A1(G78), .A2(n784), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n549), .A2(n548), .ZN(n553) );
  NAND2_X1 U607 ( .A1(n788), .A2(G53), .ZN(n551) );
  NAND2_X1 U608 ( .A1(G65), .A2(n789), .ZN(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n552) );
  OR2_X1 U610 ( .A1(n553), .A2(n552), .ZN(G299) );
  NAND2_X1 U611 ( .A1(G64), .A2(n789), .ZN(n554) );
  XNOR2_X1 U612 ( .A(KEYINPUT67), .B(n554), .ZN(n561) );
  NAND2_X1 U613 ( .A1(G90), .A2(n783), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G77), .A2(n784), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U616 ( .A(n557), .B(KEYINPUT9), .ZN(n559) );
  NAND2_X1 U617 ( .A1(G52), .A2(n788), .ZN(n558) );
  NAND2_X1 U618 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U619 ( .A1(n561), .A2(n560), .ZN(G171) );
  INV_X1 U620 ( .A(G171), .ZN(G301) );
  NAND2_X1 U621 ( .A1(n788), .A2(G51), .ZN(n563) );
  NAND2_X1 U622 ( .A1(G63), .A2(n789), .ZN(n562) );
  NAND2_X1 U623 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U624 ( .A(KEYINPUT6), .B(n564), .ZN(n571) );
  NAND2_X1 U625 ( .A1(n783), .A2(G89), .ZN(n565) );
  XNOR2_X1 U626 ( .A(n565), .B(KEYINPUT4), .ZN(n567) );
  NAND2_X1 U627 ( .A1(G76), .A2(n784), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U629 ( .A(KEYINPUT73), .B(n568), .ZN(n569) );
  XNOR2_X1 U630 ( .A(KEYINPUT5), .B(n569), .ZN(n570) );
  NOR2_X1 U631 ( .A1(n571), .A2(n570), .ZN(n572) );
  XOR2_X1 U632 ( .A(KEYINPUT7), .B(n572), .Z(G168) );
  NAND2_X1 U633 ( .A1(G88), .A2(n783), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G75), .A2(n784), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U636 ( .A(KEYINPUT81), .B(n575), .ZN(n579) );
  NAND2_X1 U637 ( .A1(n789), .A2(G62), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n788), .A2(G50), .ZN(n576) );
  AND2_X1 U639 ( .A1(n577), .A2(n576), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n579), .A2(n578), .ZN(G303) );
  XOR2_X1 U641 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U642 ( .A1(G85), .A2(n783), .ZN(n581) );
  NAND2_X1 U643 ( .A1(G60), .A2(n789), .ZN(n580) );
  NAND2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U645 ( .A1(G72), .A2(n784), .ZN(n582) );
  XNOR2_X1 U646 ( .A(KEYINPUT65), .B(n582), .ZN(n583) );
  NOR2_X1 U647 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U648 ( .A1(n788), .A2(G47), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n586), .A2(n585), .ZN(G290) );
  XOR2_X1 U650 ( .A(G1981), .B(G305), .Z(n917) );
  NOR2_X2 U651 ( .A1(G164), .A2(G1384), .ZN(n709) );
  NAND2_X1 U652 ( .A1(G160), .A2(G40), .ZN(n710) );
  INV_X1 U653 ( .A(n710), .ZN(n587) );
  NAND2_X2 U654 ( .A1(n709), .A2(n587), .ZN(n649) );
  NAND2_X1 U655 ( .A1(G8), .A2(n649), .ZN(n689) );
  NOR2_X1 U656 ( .A1(G1976), .A2(G288), .ZN(n673) );
  NAND2_X1 U657 ( .A1(n673), .A2(KEYINPUT33), .ZN(n588) );
  NOR2_X1 U658 ( .A1(n689), .A2(n588), .ZN(n678) );
  NAND2_X1 U659 ( .A1(G79), .A2(n784), .ZN(n590) );
  NAND2_X1 U660 ( .A1(G54), .A2(n788), .ZN(n589) );
  NAND2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G92), .A2(n783), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G66), .A2(n789), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n593) );
  XOR2_X1 U665 ( .A(KEYINPUT71), .B(n593), .Z(n594) );
  NOR2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X2 U667 ( .A(KEYINPUT15), .B(n596), .Z(n913) );
  NAND2_X1 U668 ( .A1(n783), .A2(G81), .ZN(n597) );
  XNOR2_X1 U669 ( .A(KEYINPUT12), .B(n597), .ZN(n600) );
  NAND2_X1 U670 ( .A1(n784), .A2(G68), .ZN(n598) );
  XOR2_X1 U671 ( .A(KEYINPUT69), .B(n598), .Z(n599) );
  NAND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n601) );
  XNOR2_X1 U673 ( .A(KEYINPUT13), .B(n601), .ZN(n607) );
  NAND2_X1 U674 ( .A1(n789), .A2(G56), .ZN(n602) );
  XOR2_X1 U675 ( .A(KEYINPUT14), .B(n602), .Z(n605) );
  NAND2_X1 U676 ( .A1(n788), .A2(G43), .ZN(n603) );
  XOR2_X1 U677 ( .A(KEYINPUT70), .B(n603), .Z(n604) );
  NOR2_X1 U678 ( .A1(n605), .A2(n604), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n607), .A2(n606), .ZN(n914) );
  INV_X1 U680 ( .A(G1996), .ZN(n727) );
  NOR2_X1 U681 ( .A1(n649), .A2(n727), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n609), .B(n608), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n649), .A2(G1341), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U685 ( .A1(n914), .A2(n612), .ZN(n618) );
  NAND2_X1 U686 ( .A1(n913), .A2(n618), .ZN(n617) );
  NAND2_X1 U687 ( .A1(G1348), .A2(n649), .ZN(n615) );
  INV_X1 U688 ( .A(n649), .ZN(n634) );
  NAND2_X1 U689 ( .A1(G2067), .A2(n623), .ZN(n614) );
  NAND2_X1 U690 ( .A1(n615), .A2(n614), .ZN(n616) );
  AND2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n620) );
  NOR2_X1 U692 ( .A1(n913), .A2(n618), .ZN(n619) );
  NOR2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n627) );
  XNOR2_X1 U694 ( .A(KEYINPUT27), .B(KEYINPUT92), .ZN(n621) );
  XNOR2_X1 U695 ( .A(n622), .B(n621), .ZN(n625) );
  INV_X1 U696 ( .A(n623), .ZN(n636) );
  NAND2_X1 U697 ( .A1(n636), .A2(G1956), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n625), .A2(n624), .ZN(n629) );
  NOR2_X1 U699 ( .A1(G299), .A2(n629), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U701 ( .A(KEYINPUT93), .B(n628), .Z(n632) );
  NAND2_X1 U702 ( .A1(G299), .A2(n629), .ZN(n630) );
  XOR2_X1 U703 ( .A(KEYINPUT28), .B(n630), .Z(n631) );
  XNOR2_X1 U704 ( .A(n633), .B(KEYINPUT29), .ZN(n640) );
  NOR2_X1 U705 ( .A1(n634), .A2(G1961), .ZN(n635) );
  XNOR2_X1 U706 ( .A(n635), .B(KEYINPUT90), .ZN(n638) );
  XOR2_X1 U707 ( .A(G2078), .B(KEYINPUT25), .Z(n970) );
  NOR2_X1 U708 ( .A1(n636), .A2(n970), .ZN(n637) );
  NOR2_X1 U709 ( .A1(n638), .A2(n637), .ZN(n645) );
  OR2_X1 U710 ( .A1(G301), .A2(n645), .ZN(n639) );
  NAND2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n664) );
  NOR2_X1 U712 ( .A1(G1966), .A2(n689), .ZN(n666) );
  NOR2_X1 U713 ( .A1(G2084), .A2(n649), .ZN(n662) );
  NOR2_X1 U714 ( .A1(n666), .A2(n662), .ZN(n641) );
  NAND2_X1 U715 ( .A1(G8), .A2(n641), .ZN(n642) );
  XNOR2_X1 U716 ( .A(KEYINPUT30), .B(n642), .ZN(n643) );
  NOR2_X1 U717 ( .A1(G168), .A2(n643), .ZN(n644) );
  XOR2_X1 U718 ( .A(KEYINPUT94), .B(n644), .Z(n647) );
  NAND2_X1 U719 ( .A1(n645), .A2(G301), .ZN(n646) );
  NAND2_X1 U720 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n648), .B(KEYINPUT31), .ZN(n665) );
  INV_X1 U722 ( .A(G8), .ZN(n654) );
  NOR2_X1 U723 ( .A1(G1971), .A2(n689), .ZN(n651) );
  NOR2_X1 U724 ( .A1(G2090), .A2(n649), .ZN(n650) );
  NOR2_X1 U725 ( .A1(n651), .A2(n650), .ZN(n652) );
  NAND2_X1 U726 ( .A1(n652), .A2(G303), .ZN(n653) );
  OR2_X1 U727 ( .A1(n654), .A2(n653), .ZN(n656) );
  AND2_X1 U728 ( .A1(n665), .A2(n656), .ZN(n655) );
  NAND2_X1 U729 ( .A1(n664), .A2(n655), .ZN(n660) );
  INV_X1 U730 ( .A(n656), .ZN(n658) );
  AND2_X1 U731 ( .A1(G286), .A2(G8), .ZN(n657) );
  OR2_X1 U732 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U734 ( .A1(G8), .A2(n662), .ZN(n663) );
  XOR2_X1 U735 ( .A(KEYINPUT89), .B(n663), .Z(n669) );
  AND2_X1 U736 ( .A1(n665), .A2(n664), .ZN(n667) );
  NOR2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U738 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n687) );
  NOR2_X1 U740 ( .A1(G1971), .A2(G303), .ZN(n672) );
  NOR2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n930) );
  NAND2_X1 U742 ( .A1(n687), .A2(n930), .ZN(n674) );
  NAND2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n924) );
  NAND2_X1 U744 ( .A1(n674), .A2(n924), .ZN(n675) );
  NOR2_X1 U745 ( .A1(KEYINPUT33), .A2(n676), .ZN(n677) );
  NOR2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n679) );
  NAND2_X1 U747 ( .A1(n917), .A2(n679), .ZN(n680) );
  XNOR2_X1 U748 ( .A(n680), .B(KEYINPUT95), .ZN(n684) );
  NOR2_X1 U749 ( .A1(G1981), .A2(G305), .ZN(n681) );
  XOR2_X1 U750 ( .A(n681), .B(KEYINPUT24), .Z(n682) );
  NOR2_X1 U751 ( .A1(n689), .A2(n682), .ZN(n683) );
  NOR2_X1 U752 ( .A1(G2090), .A2(G303), .ZN(n685) );
  NAND2_X1 U753 ( .A1(G8), .A2(n685), .ZN(n686) );
  NAND2_X1 U754 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n690) );
  NAND2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n725) );
  XOR2_X1 U757 ( .A(G1986), .B(G290), .Z(n926) );
  XOR2_X1 U758 ( .A(KEYINPUT86), .B(G1991), .Z(n967) );
  NAND2_X1 U759 ( .A1(G131), .A2(n885), .ZN(n693) );
  NAND2_X1 U760 ( .A1(G95), .A2(n883), .ZN(n692) );
  NAND2_X1 U761 ( .A1(n693), .A2(n692), .ZN(n697) );
  NAND2_X1 U762 ( .A1(G107), .A2(n879), .ZN(n695) );
  NAND2_X1 U763 ( .A1(G119), .A2(n880), .ZN(n694) );
  NAND2_X1 U764 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U765 ( .A1(n697), .A2(n696), .ZN(n876) );
  NOR2_X1 U766 ( .A1(n967), .A2(n876), .ZN(n698) );
  XOR2_X1 U767 ( .A(KEYINPUT87), .B(n698), .Z(n708) );
  NAND2_X1 U768 ( .A1(G105), .A2(n883), .ZN(n699) );
  XNOR2_X1 U769 ( .A(n699), .B(KEYINPUT38), .ZN(n700) );
  XNOR2_X1 U770 ( .A(n700), .B(KEYINPUT88), .ZN(n702) );
  NAND2_X1 U771 ( .A1(G117), .A2(n879), .ZN(n701) );
  NAND2_X1 U772 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U773 ( .A1(G141), .A2(n885), .ZN(n704) );
  NAND2_X1 U774 ( .A1(G129), .A2(n880), .ZN(n703) );
  NAND2_X1 U775 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U776 ( .A1(n706), .A2(n705), .ZN(n891) );
  NOR2_X1 U777 ( .A1(n891), .A2(n727), .ZN(n707) );
  NOR2_X1 U778 ( .A1(n708), .A2(n707), .ZN(n992) );
  NAND2_X1 U779 ( .A1(n926), .A2(n992), .ZN(n711) );
  NOR2_X1 U780 ( .A1(n710), .A2(n709), .ZN(n740) );
  NAND2_X1 U781 ( .A1(n711), .A2(n740), .ZN(n723) );
  XOR2_X1 U782 ( .A(KEYINPUT37), .B(G2067), .Z(n739) );
  NAND2_X1 U783 ( .A1(n885), .A2(G140), .ZN(n712) );
  XNOR2_X1 U784 ( .A(n712), .B(KEYINPUT84), .ZN(n714) );
  NAND2_X1 U785 ( .A1(G104), .A2(n883), .ZN(n713) );
  NAND2_X1 U786 ( .A1(n714), .A2(n713), .ZN(n715) );
  XNOR2_X1 U787 ( .A(KEYINPUT34), .B(n715), .ZN(n721) );
  NAND2_X1 U788 ( .A1(G116), .A2(n879), .ZN(n717) );
  NAND2_X1 U789 ( .A1(G128), .A2(n880), .ZN(n716) );
  NAND2_X1 U790 ( .A1(n717), .A2(n716), .ZN(n718) );
  XNOR2_X1 U791 ( .A(KEYINPUT85), .B(n718), .ZN(n719) );
  XNOR2_X1 U792 ( .A(KEYINPUT35), .B(n719), .ZN(n720) );
  NOR2_X1 U793 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U794 ( .A(KEYINPUT36), .B(n722), .Z(n895) );
  AND2_X1 U795 ( .A1(n739), .A2(n895), .ZN(n990) );
  NAND2_X1 U796 ( .A1(n990), .A2(n740), .ZN(n726) );
  AND2_X1 U797 ( .A1(n723), .A2(n726), .ZN(n724) );
  NAND2_X1 U798 ( .A1(n725), .A2(n724), .ZN(n738) );
  INV_X1 U799 ( .A(n726), .ZN(n736) );
  AND2_X1 U800 ( .A1(n727), .A2(n891), .ZN(n987) );
  NOR2_X1 U801 ( .A1(G1986), .A2(G290), .ZN(n729) );
  NAND2_X1 U802 ( .A1(n876), .A2(n967), .ZN(n728) );
  XOR2_X1 U803 ( .A(KEYINPUT96), .B(n728), .Z(n993) );
  NOR2_X1 U804 ( .A1(n729), .A2(n993), .ZN(n731) );
  INV_X1 U805 ( .A(n992), .ZN(n730) );
  NOR2_X1 U806 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U807 ( .A1(n987), .A2(n732), .ZN(n733) );
  XNOR2_X1 U808 ( .A(KEYINPUT39), .B(n733), .ZN(n734) );
  NAND2_X1 U809 ( .A1(n734), .A2(n740), .ZN(n735) );
  OR2_X1 U810 ( .A1(n736), .A2(n735), .ZN(n737) );
  AND2_X1 U811 ( .A1(n738), .A2(n737), .ZN(n742) );
  NOR2_X1 U812 ( .A1(n739), .A2(n895), .ZN(n1005) );
  NAND2_X1 U813 ( .A1(n1005), .A2(n740), .ZN(n741) );
  NAND2_X1 U814 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U815 ( .A(n743), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U816 ( .A(G2451), .B(G2427), .ZN(n753) );
  XOR2_X1 U817 ( .A(G2430), .B(G2443), .Z(n745) );
  XNOR2_X1 U818 ( .A(G2435), .B(G2438), .ZN(n744) );
  XNOR2_X1 U819 ( .A(n745), .B(n744), .ZN(n749) );
  XOR2_X1 U820 ( .A(G2454), .B(KEYINPUT97), .Z(n747) );
  XNOR2_X1 U821 ( .A(G1341), .B(G1348), .ZN(n746) );
  XNOR2_X1 U822 ( .A(n747), .B(n746), .ZN(n748) );
  XOR2_X1 U823 ( .A(n749), .B(n748), .Z(n751) );
  XNOR2_X1 U824 ( .A(G2446), .B(KEYINPUT98), .ZN(n750) );
  XNOR2_X1 U825 ( .A(n751), .B(n750), .ZN(n752) );
  XNOR2_X1 U826 ( .A(n753), .B(n752), .ZN(n754) );
  AND2_X1 U827 ( .A1(n754), .A2(G14), .ZN(G401) );
  AND2_X1 U828 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U829 ( .A(G108), .ZN(G238) );
  INV_X1 U830 ( .A(G69), .ZN(G235) );
  INV_X1 U831 ( .A(G132), .ZN(G219) );
  INV_X1 U832 ( .A(G82), .ZN(G220) );
  NAND2_X1 U833 ( .A1(G7), .A2(G661), .ZN(n755) );
  XNOR2_X1 U834 ( .A(n755), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U835 ( .A(G567), .ZN(n818) );
  NOR2_X1 U836 ( .A1(n818), .A2(G223), .ZN(n756) );
  XNOR2_X1 U837 ( .A(n756), .B(KEYINPUT11), .ZN(G234) );
  INV_X1 U838 ( .A(G860), .ZN(n765) );
  OR2_X1 U839 ( .A1(n914), .A2(n765), .ZN(G153) );
  NOR2_X1 U840 ( .A1(n913), .A2(G868), .ZN(n757) );
  XOR2_X1 U841 ( .A(KEYINPUT72), .B(n757), .Z(n759) );
  NAND2_X1 U842 ( .A1(G868), .A2(G301), .ZN(n758) );
  NAND2_X1 U843 ( .A1(n759), .A2(n758), .ZN(G284) );
  INV_X1 U844 ( .A(G868), .ZN(n803) );
  XNOR2_X1 U845 ( .A(KEYINPUT74), .B(n803), .ZN(n760) );
  NOR2_X1 U846 ( .A1(G286), .A2(n760), .ZN(n761) );
  XOR2_X1 U847 ( .A(KEYINPUT75), .B(n761), .Z(n764) );
  NOR2_X1 U848 ( .A1(G868), .A2(G299), .ZN(n762) );
  XNOR2_X1 U849 ( .A(KEYINPUT76), .B(n762), .ZN(n763) );
  NOR2_X1 U850 ( .A1(n764), .A2(n763), .ZN(G297) );
  NAND2_X1 U851 ( .A1(n765), .A2(G559), .ZN(n766) );
  NAND2_X1 U852 ( .A1(n766), .A2(n913), .ZN(n767) );
  XNOR2_X1 U853 ( .A(n767), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U854 ( .A1(G868), .A2(n914), .ZN(n770) );
  NAND2_X1 U855 ( .A1(G868), .A2(n913), .ZN(n768) );
  NOR2_X1 U856 ( .A1(G559), .A2(n768), .ZN(n769) );
  NOR2_X1 U857 ( .A1(n770), .A2(n769), .ZN(G282) );
  NAND2_X1 U858 ( .A1(G99), .A2(n883), .ZN(n772) );
  NAND2_X1 U859 ( .A1(G111), .A2(n879), .ZN(n771) );
  NAND2_X1 U860 ( .A1(n772), .A2(n771), .ZN(n779) );
  NAND2_X1 U861 ( .A1(n885), .A2(G135), .ZN(n773) );
  XNOR2_X1 U862 ( .A(KEYINPUT77), .B(n773), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n880), .A2(G123), .ZN(n774) );
  XOR2_X1 U864 ( .A(KEYINPUT18), .B(n774), .Z(n775) );
  NOR2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U866 ( .A(KEYINPUT78), .B(n777), .Z(n778) );
  NOR2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n994) );
  XNOR2_X1 U868 ( .A(n994), .B(G2096), .ZN(n781) );
  INV_X1 U869 ( .A(G2100), .ZN(n780) );
  NAND2_X1 U870 ( .A1(n781), .A2(n780), .ZN(G156) );
  NAND2_X1 U871 ( .A1(n913), .A2(G559), .ZN(n801) );
  XNOR2_X1 U872 ( .A(n914), .B(n801), .ZN(n782) );
  NOR2_X1 U873 ( .A1(n782), .A2(G860), .ZN(n794) );
  NAND2_X1 U874 ( .A1(n783), .A2(G93), .ZN(n787) );
  NAND2_X1 U875 ( .A1(G80), .A2(n784), .ZN(n785) );
  XOR2_X1 U876 ( .A(KEYINPUT79), .B(n785), .Z(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n793) );
  NAND2_X1 U878 ( .A1(n788), .A2(G55), .ZN(n791) );
  NAND2_X1 U879 ( .A1(G67), .A2(n789), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n792) );
  OR2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n804) );
  XOR2_X1 U882 ( .A(n794), .B(n804), .Z(G145) );
  INV_X1 U883 ( .A(G303), .ZN(G166) );
  XNOR2_X1 U884 ( .A(G166), .B(G299), .ZN(n795) );
  XNOR2_X1 U885 ( .A(n795), .B(G290), .ZN(n796) );
  XNOR2_X1 U886 ( .A(n796), .B(n914), .ZN(n797) );
  XNOR2_X1 U887 ( .A(n797), .B(G305), .ZN(n798) );
  XOR2_X1 U888 ( .A(n804), .B(n798), .Z(n800) );
  XNOR2_X1 U889 ( .A(G288), .B(KEYINPUT19), .ZN(n799) );
  XNOR2_X1 U890 ( .A(n800), .B(n799), .ZN(n899) );
  XOR2_X1 U891 ( .A(n899), .B(n801), .Z(n802) );
  NAND2_X1 U892 ( .A1(G868), .A2(n802), .ZN(n806) );
  NAND2_X1 U893 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U894 ( .A1(n806), .A2(n805), .ZN(G295) );
  NAND2_X1 U895 ( .A1(G2078), .A2(G2084), .ZN(n807) );
  XOR2_X1 U896 ( .A(KEYINPUT20), .B(n807), .Z(n808) );
  NAND2_X1 U897 ( .A1(G2090), .A2(n808), .ZN(n809) );
  XNOR2_X1 U898 ( .A(KEYINPUT21), .B(n809), .ZN(n810) );
  NAND2_X1 U899 ( .A1(n810), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U900 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U901 ( .A(KEYINPUT68), .B(G57), .Z(G237) );
  NOR2_X1 U902 ( .A1(G220), .A2(G219), .ZN(n811) );
  XOR2_X1 U903 ( .A(KEYINPUT22), .B(n811), .Z(n812) );
  NOR2_X1 U904 ( .A1(G218), .A2(n812), .ZN(n813) );
  XNOR2_X1 U905 ( .A(KEYINPUT82), .B(n813), .ZN(n814) );
  NAND2_X1 U906 ( .A1(n814), .A2(G96), .ZN(n829) );
  NAND2_X1 U907 ( .A1(G2106), .A2(n829), .ZN(n815) );
  XNOR2_X1 U908 ( .A(n815), .B(KEYINPUT83), .ZN(n820) );
  NOR2_X1 U909 ( .A1(G237), .A2(G238), .ZN(n816) );
  NAND2_X1 U910 ( .A1(G120), .A2(n816), .ZN(n817) );
  NOR2_X1 U911 ( .A1(G235), .A2(n817), .ZN(n828) );
  NOR2_X1 U912 ( .A1(n818), .A2(n828), .ZN(n819) );
  NOR2_X1 U913 ( .A1(n820), .A2(n819), .ZN(G319) );
  INV_X1 U914 ( .A(G319), .ZN(n822) );
  NAND2_X1 U915 ( .A1(G483), .A2(G661), .ZN(n821) );
  NOR2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n827) );
  NAND2_X1 U917 ( .A1(n827), .A2(G36), .ZN(G176) );
  INV_X1 U918 ( .A(G223), .ZN(n823) );
  NAND2_X1 U919 ( .A1(n823), .A2(G2106), .ZN(n824) );
  XOR2_X1 U920 ( .A(KEYINPUT99), .B(n824), .Z(G217) );
  AND2_X1 U921 ( .A1(G15), .A2(G2), .ZN(n825) );
  NAND2_X1 U922 ( .A1(G661), .A2(n825), .ZN(G259) );
  NAND2_X1 U923 ( .A1(G3), .A2(G1), .ZN(n826) );
  NAND2_X1 U924 ( .A1(n827), .A2(n826), .ZN(G188) );
  INV_X1 U925 ( .A(n828), .ZN(n830) );
  NOR2_X1 U926 ( .A1(n830), .A2(n829), .ZN(G325) );
  XOR2_X1 U927 ( .A(KEYINPUT100), .B(G325), .Z(G261) );
  INV_X1 U929 ( .A(G96), .ZN(G221) );
  XOR2_X1 U930 ( .A(KEYINPUT42), .B(G2090), .Z(n832) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2084), .ZN(n831) );
  XNOR2_X1 U932 ( .A(n832), .B(n831), .ZN(n833) );
  XOR2_X1 U933 ( .A(n833), .B(G2100), .Z(n835) );
  XNOR2_X1 U934 ( .A(G2078), .B(G2072), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n835), .B(n834), .ZN(n839) );
  XOR2_X1 U936 ( .A(G2096), .B(KEYINPUT43), .Z(n837) );
  XNOR2_X1 U937 ( .A(G2678), .B(KEYINPUT101), .ZN(n836) );
  XNOR2_X1 U938 ( .A(n837), .B(n836), .ZN(n838) );
  XOR2_X1 U939 ( .A(n839), .B(n838), .Z(G227) );
  XOR2_X1 U940 ( .A(KEYINPUT102), .B(KEYINPUT41), .Z(n841) );
  XNOR2_X1 U941 ( .A(KEYINPUT103), .B(KEYINPUT104), .ZN(n840) );
  XNOR2_X1 U942 ( .A(n841), .B(n840), .ZN(n842) );
  XOR2_X1 U943 ( .A(n842), .B(G2474), .Z(n844) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1981), .ZN(n843) );
  XNOR2_X1 U945 ( .A(n844), .B(n843), .ZN(n852) );
  XOR2_X1 U946 ( .A(G1986), .B(G1976), .Z(n846) );
  XNOR2_X1 U947 ( .A(G1956), .B(G1971), .ZN(n845) );
  XNOR2_X1 U948 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U949 ( .A(KEYINPUT105), .B(G1991), .Z(n848) );
  XNOR2_X1 U950 ( .A(G1961), .B(G1996), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U952 ( .A(n850), .B(n849), .Z(n851) );
  XNOR2_X1 U953 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U954 ( .A1(G124), .A2(n880), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n853), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U956 ( .A1(G100), .A2(n883), .ZN(n854) );
  XNOR2_X1 U957 ( .A(n854), .B(KEYINPUT106), .ZN(n855) );
  NAND2_X1 U958 ( .A1(n856), .A2(n855), .ZN(n860) );
  NAND2_X1 U959 ( .A1(G136), .A2(n885), .ZN(n858) );
  NAND2_X1 U960 ( .A1(G112), .A2(n879), .ZN(n857) );
  NAND2_X1 U961 ( .A1(n858), .A2(n857), .ZN(n859) );
  NOR2_X1 U962 ( .A1(n860), .A2(n859), .ZN(G162) );
  XOR2_X1 U963 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n862) );
  XNOR2_X1 U964 ( .A(G164), .B(n994), .ZN(n861) );
  XNOR2_X1 U965 ( .A(n862), .B(n861), .ZN(n875) );
  NAND2_X1 U966 ( .A1(n880), .A2(G127), .ZN(n863) );
  XNOR2_X1 U967 ( .A(KEYINPUT110), .B(n863), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n879), .A2(G115), .ZN(n864) );
  XOR2_X1 U969 ( .A(KEYINPUT111), .B(n864), .Z(n865) );
  NAND2_X1 U970 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U971 ( .A(n867), .B(KEYINPUT47), .ZN(n873) );
  NAND2_X1 U972 ( .A1(n885), .A2(G139), .ZN(n868) );
  XNOR2_X1 U973 ( .A(n868), .B(KEYINPUT108), .ZN(n870) );
  NAND2_X1 U974 ( .A1(G103), .A2(n883), .ZN(n869) );
  NAND2_X1 U975 ( .A1(n870), .A2(n869), .ZN(n871) );
  XNOR2_X1 U976 ( .A(KEYINPUT109), .B(n871), .ZN(n872) );
  NAND2_X1 U977 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U978 ( .A(n874), .B(KEYINPUT112), .ZN(n1000) );
  XOR2_X1 U979 ( .A(n875), .B(n1000), .Z(n878) );
  XNOR2_X1 U980 ( .A(G160), .B(n876), .ZN(n877) );
  XNOR2_X1 U981 ( .A(n878), .B(n877), .ZN(n894) );
  NAND2_X1 U982 ( .A1(G118), .A2(n879), .ZN(n882) );
  NAND2_X1 U983 ( .A1(G130), .A2(n880), .ZN(n881) );
  NAND2_X1 U984 ( .A1(n882), .A2(n881), .ZN(n890) );
  NAND2_X1 U985 ( .A1(n883), .A2(G106), .ZN(n884) );
  XOR2_X1 U986 ( .A(KEYINPUT107), .B(n884), .Z(n887) );
  NAND2_X1 U987 ( .A1(n885), .A2(G142), .ZN(n886) );
  NAND2_X1 U988 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U989 ( .A(n888), .B(KEYINPUT45), .Z(n889) );
  NOR2_X1 U990 ( .A1(n890), .A2(n889), .ZN(n892) );
  XOR2_X1 U991 ( .A(n892), .B(n891), .Z(n893) );
  XOR2_X1 U992 ( .A(n894), .B(n893), .Z(n897) );
  XNOR2_X1 U993 ( .A(n895), .B(G162), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n898) );
  NOR2_X1 U995 ( .A1(G37), .A2(n898), .ZN(G395) );
  XOR2_X1 U996 ( .A(KEYINPUT113), .B(n899), .Z(n901) );
  XNOR2_X1 U997 ( .A(G171), .B(G286), .ZN(n900) );
  XNOR2_X1 U998 ( .A(n901), .B(n900), .ZN(n902) );
  XNOR2_X1 U999 ( .A(n902), .B(n913), .ZN(n903) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n903), .ZN(G397) );
  NOR2_X1 U1001 ( .A1(G227), .A2(G229), .ZN(n904) );
  XOR2_X1 U1002 ( .A(KEYINPUT49), .B(n904), .Z(n905) );
  NAND2_X1 U1003 ( .A1(G319), .A2(n905), .ZN(n906) );
  NOR2_X1 U1004 ( .A1(G401), .A2(n906), .ZN(n907) );
  XOR2_X1 U1005 ( .A(KEYINPUT114), .B(n907), .Z(n910) );
  NOR2_X1 U1006 ( .A1(G395), .A2(G397), .ZN(n908) );
  XNOR2_X1 U1007 ( .A(KEYINPUT115), .B(n908), .ZN(n909) );
  NOR2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(KEYINPUT116), .B(n911), .ZN(G308) );
  INV_X1 U1010 ( .A(G308), .ZN(G225) );
  INV_X1 U1011 ( .A(G120), .ZN(G236) );
  XNOR2_X1 U1012 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n1017) );
  XNOR2_X1 U1013 ( .A(G16), .B(KEYINPUT122), .ZN(n912) );
  XNOR2_X1 U1014 ( .A(n912), .B(KEYINPUT56), .ZN(n936) );
  XNOR2_X1 U1015 ( .A(n913), .B(G1348), .ZN(n916) );
  XOR2_X1 U1016 ( .A(G1341), .B(n914), .Z(n915) );
  NAND2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n922) );
  XNOR2_X1 U1018 ( .A(G1966), .B(G168), .ZN(n918) );
  NAND2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(n919), .B(KEYINPUT57), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(n920), .B(KEYINPUT123), .ZN(n921) );
  NOR2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n934) );
  XOR2_X1 U1023 ( .A(G1956), .B(G299), .Z(n923) );
  NAND2_X1 U1024 ( .A1(n924), .A2(n923), .ZN(n932) );
  NAND2_X1 U1025 ( .A1(G1971), .A2(G303), .ZN(n925) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n928) );
  XNOR2_X1 U1027 ( .A(G1961), .B(G301), .ZN(n927) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1030 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1031 ( .A1(n934), .A2(n933), .ZN(n935) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1033 ( .A(KEYINPUT124), .B(n937), .ZN(n1015) );
  XNOR2_X1 U1034 ( .A(G1971), .B(G22), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(G23), .B(G1976), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n941) );
  XOR2_X1 U1037 ( .A(G1986), .B(G24), .Z(n940) );
  NAND2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n943) );
  XOR2_X1 U1039 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n942) );
  XNOR2_X1 U1040 ( .A(n943), .B(n942), .ZN(n956) );
  XNOR2_X1 U1041 ( .A(G1348), .B(KEYINPUT59), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(n944), .B(G4), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(G1956), .B(G20), .ZN(n946) );
  XNOR2_X1 U1044 ( .A(G6), .B(G1981), .ZN(n945) );
  NOR2_X1 U1045 ( .A1(n946), .A2(n945), .ZN(n947) );
  NAND2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n951) );
  XOR2_X1 U1047 ( .A(KEYINPUT125), .B(G1341), .Z(n949) );
  XNOR2_X1 U1048 ( .A(G19), .B(n949), .ZN(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  XOR2_X1 U1050 ( .A(KEYINPUT60), .B(n952), .Z(n954) );
  XNOR2_X1 U1051 ( .A(G1966), .B(G21), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n958) );
  XNOR2_X1 U1054 ( .A(G5), .B(G1961), .ZN(n957) );
  NOR2_X1 U1055 ( .A1(n958), .A2(n957), .ZN(n959) );
  XNOR2_X1 U1056 ( .A(KEYINPUT61), .B(n959), .ZN(n961) );
  INV_X1 U1057 ( .A(G16), .ZN(n960) );
  NAND2_X1 U1058 ( .A1(n961), .A2(n960), .ZN(n962) );
  NAND2_X1 U1059 ( .A1(n962), .A2(G11), .ZN(n1013) );
  XOR2_X1 U1060 ( .A(G2090), .B(G35), .Z(n980) );
  XNOR2_X1 U1061 ( .A(G2072), .B(G33), .ZN(n963) );
  XNOR2_X1 U1062 ( .A(n963), .B(KEYINPUT118), .ZN(n965) );
  XNOR2_X1 U1063 ( .A(G26), .B(G2067), .ZN(n964) );
  NOR2_X1 U1064 ( .A1(n965), .A2(n964), .ZN(n966) );
  XOR2_X1 U1065 ( .A(KEYINPUT119), .B(n966), .Z(n969) );
  XNOR2_X1 U1066 ( .A(n967), .B(G25), .ZN(n968) );
  NAND2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n970), .B(G27), .ZN(n972) );
  XNOR2_X1 U1069 ( .A(G32), .B(G1996), .ZN(n971) );
  NOR2_X1 U1070 ( .A1(n972), .A2(n971), .ZN(n973) );
  XOR2_X1 U1071 ( .A(KEYINPUT120), .B(n973), .Z(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1073 ( .A1(n976), .A2(G28), .ZN(n977) );
  XOR2_X1 U1074 ( .A(KEYINPUT53), .B(n977), .Z(n978) );
  XNOR2_X1 U1075 ( .A(n978), .B(KEYINPUT121), .ZN(n979) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n983) );
  XNOR2_X1 U1077 ( .A(G34), .B(G2084), .ZN(n981) );
  XNOR2_X1 U1078 ( .A(KEYINPUT54), .B(n981), .ZN(n982) );
  NOR2_X1 U1079 ( .A1(n983), .A2(n982), .ZN(n984) );
  NOR2_X1 U1080 ( .A1(G29), .A2(n984), .ZN(n985) );
  XNOR2_X1 U1081 ( .A(n985), .B(KEYINPUT55), .ZN(n1011) );
  XOR2_X1 U1082 ( .A(G2090), .B(G162), .Z(n986) );
  NOR2_X1 U1083 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1084 ( .A(n988), .B(KEYINPUT51), .ZN(n989) );
  NOR2_X1 U1085 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n999) );
  NOR2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(G160), .B(G2084), .ZN(n995) );
  NAND2_X1 U1089 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1090 ( .A(KEYINPUT117), .B(n997), .Z(n998) );
  NOR2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1007) );
  XOR2_X1 U1092 ( .A(G164), .B(G2078), .Z(n1002) );
  XNOR2_X1 U1093 ( .A(G2072), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1095 ( .A(KEYINPUT50), .B(n1003), .Z(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1097 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  XNOR2_X1 U1098 ( .A(KEYINPUT52), .B(n1008), .ZN(n1009) );
  NAND2_X1 U1099 ( .A1(G29), .A2(n1009), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(n1017), .B(n1016), .ZN(G311) );
  INV_X1 U1104 ( .A(G311), .ZN(G150) );
endmodule

