//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:43 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n564, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n573, new_n574, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT64), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(KEYINPUT65), .B(KEYINPUT2), .Z(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n453), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(KEYINPUT67), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n462), .B1(KEYINPUT3), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g039(.A(KEYINPUT66), .B(KEYINPUT3), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n464), .B1(new_n465), .B2(new_n463), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT3), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n469), .A2(KEYINPUT66), .ZN(new_n470));
  OAI211_X1 g045(.A(new_n462), .B(G2104), .C1(new_n468), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  XNOR2_X1  g051(.A(KEYINPUT3), .B(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G125), .ZN(new_n478));
  INV_X1    g053(.A(G113), .ZN(new_n479));
  OAI21_X1  g054(.A(new_n478), .B1(new_n479), .B2(new_n463), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n463), .A2(G2105), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n480), .A2(G2105), .B1(G101), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G160));
  NAND2_X1  g059(.A1(new_n475), .A2(G136), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n472), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n473), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NAND4_X1  g067(.A1(new_n472), .A2(KEYINPUT4), .A3(G138), .A4(new_n473), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n477), .A2(G138), .A3(new_n473), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  INV_X1    g073(.A(G114), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(G126), .A2(G2105), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g078(.A(KEYINPUT68), .B1(new_n472), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT68), .ZN(new_n505));
  AOI211_X1 g080(.A(new_n505), .B(new_n502), .C1(new_n466), .C2(new_n471), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT69), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g084(.A(KEYINPUT69), .B(new_n501), .C1(new_n504), .C2(new_n506), .ZN(new_n510));
  AOI21_X1  g085(.A(new_n497), .B1(new_n509), .B2(new_n510), .ZN(G164));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT6), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT70), .A2(KEYINPUT6), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n512), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT71), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(KEYINPUT71), .B1(new_n514), .B2(G651), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n521), .A2(G543), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n524));
  INV_X1    g099(.A(G543), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n525), .B2(KEYINPUT5), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT5), .ZN(new_n527));
  NAND3_X1  g102(.A1(new_n527), .A2(KEYINPUT72), .A3(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n525), .A2(KEYINPUT5), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G62), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n523), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n522), .A2(G50), .B1(G651), .B2(new_n533), .ZN(new_n534));
  AND2_X1   g109(.A1(new_n529), .A2(new_n530), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n521), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT73), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n521), .A2(KEYINPUT73), .A3(new_n535), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(G88), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n534), .B1(new_n540), .B2(new_n541), .ZN(G303));
  INV_X1    g117(.A(G303), .ZN(G166));
  NAND3_X1  g118(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n544));
  XOR2_X1   g119(.A(new_n544), .B(KEYINPUT7), .Z(new_n545));
  AOI21_X1  g120(.A(new_n545), .B1(new_n522), .B2(G51), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT74), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n531), .B(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n548), .A2(G63), .A3(G651), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  AND3_X1   g125(.A1(new_n538), .A2(G89), .A3(new_n539), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT75), .ZN(new_n552));
  OR3_X1    g127(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n550), .B2(new_n551), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(G168));
  AND2_X1   g130(.A1(new_n538), .A2(new_n539), .ZN(new_n556));
  XOR2_X1   g131(.A(KEYINPUT76), .B(G90), .Z(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  AND2_X1   g133(.A1(new_n548), .A2(G64), .ZN(new_n559));
  AND2_X1   g134(.A1(G77), .A2(G543), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n522), .A2(G52), .ZN(new_n562));
  AND3_X1   g137(.A1(new_n558), .A2(new_n561), .A3(new_n562), .ZN(G171));
  AOI22_X1  g138(.A1(new_n556), .A2(G81), .B1(G43), .B2(new_n522), .ZN(new_n564));
  AND2_X1   g139(.A1(new_n548), .A2(G56), .ZN(new_n565));
  AND2_X1   g140(.A1(G68), .A2(G543), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(G860), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT77), .ZN(G153));
  NAND4_X1  g146(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g147(.A1(G1), .A2(G3), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT8), .ZN(new_n574));
  NAND4_X1  g149(.A1(G319), .A2(G483), .A3(G661), .A4(new_n574), .ZN(G188));
  NAND3_X1  g150(.A1(new_n521), .A2(G53), .A3(G543), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT9), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n538), .A2(G91), .A3(new_n539), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n535), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(new_n512), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  AND2_X1   g157(.A1(new_n553), .A2(new_n554), .ZN(G286));
  NAND2_X1  g158(.A1(new_n556), .A2(G87), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n522), .A2(G49), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n548), .B2(G74), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(KEYINPUT78), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n586), .A2(KEYINPUT78), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n584), .B(new_n585), .C1(new_n587), .C2(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n531), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n522), .A2(G48), .B1(G651), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(G86), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n540), .B2(new_n594), .ZN(G305));
  AOI22_X1  g170(.A1(new_n556), .A2(G85), .B1(G47), .B2(new_n522), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n548), .A2(G60), .ZN(new_n597));
  AND2_X1   g172(.A1(G72), .A2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(G651), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n596), .A2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  INV_X1    g176(.A(G54), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n521), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT79), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n604), .B2(new_n603), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n535), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n607));
  AOI21_X1  g182(.A(new_n512), .B1(new_n607), .B2(KEYINPUT80), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(KEYINPUT80), .B2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(KEYINPUT81), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n606), .A2(new_n612), .A3(new_n609), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  INV_X1    g189(.A(G92), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n540), .B2(new_n615), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n556), .A2(KEYINPUT10), .A3(G92), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n611), .A2(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n601), .B1(G868), .B2(new_n618), .ZN(G284));
  OAI21_X1  g194(.A(new_n601), .B1(G868), .B2(new_n618), .ZN(G321));
  XOR2_X1   g195(.A(G299), .B(KEYINPUT82), .Z(new_n621));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  MUX2_X1   g197(.A(G286), .B(new_n621), .S(new_n622), .Z(G280));
  XNOR2_X1  g198(.A(G280), .B(KEYINPUT83), .ZN(G297));
  XOR2_X1   g199(.A(KEYINPUT84), .B(G559), .Z(new_n625));
  OAI21_X1  g200(.A(new_n618), .B1(G860), .B2(new_n625), .ZN(G148));
  NOR2_X1   g201(.A1(new_n569), .A2(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n618), .A2(new_n625), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT85), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI211_X1 g207(.A(new_n632), .B(G2104), .C1(G111), .C2(new_n473), .ZN(new_n633));
  INV_X1    g208(.A(G135), .ZN(new_n634));
  INV_X1    g209(.A(G123), .ZN(new_n635));
  OAI221_X1 g210(.A(new_n633), .B1(new_n474), .B2(new_n634), .C1(new_n635), .C2(new_n486), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2096), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(G2096), .ZN(new_n638));
  NAND3_X1  g213(.A1(new_n473), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT12), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT13), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2100), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n637), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT86), .Z(G156));
  XNOR2_X1  g219(.A(G2427), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2430), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT15), .B(G2435), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(KEYINPUT14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1341), .B(G1348), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT87), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n650), .B(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2451), .B(G2454), .Z(new_n655));
  XNOR2_X1  g230(.A(G2443), .B(G2446), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n655), .B(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n654), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n654), .A2(new_n657), .ZN(new_n659));
  AND3_X1   g234(.A1(new_n658), .A2(G14), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT88), .Z(G401));
  INV_X1    g236(.A(KEYINPUT18), .ZN(new_n662));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(KEYINPUT17), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n663), .A2(new_n664), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n662), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(G2100), .ZN(new_n669));
  XOR2_X1   g244(.A(G2072), .B(G2078), .Z(new_n670));
  AOI21_X1  g245(.A(new_n670), .B1(new_n665), .B2(KEYINPUT18), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2096), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n669), .B(new_n672), .ZN(G227));
  XNOR2_X1  g248(.A(G1981), .B(G1986), .ZN(new_n674));
  INV_X1    g249(.A(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(G1971), .B(G1976), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT19), .ZN(new_n677));
  XOR2_X1   g252(.A(G1956), .B(G2474), .Z(new_n678));
  XOR2_X1   g253(.A(G1961), .B(G1966), .Z(new_n679));
  NOR2_X1   g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  AND2_X1   g256(.A1(new_n678), .A2(new_n679), .ZN(new_n682));
  NOR3_X1   g257(.A1(new_n677), .A2(new_n682), .A3(new_n680), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n677), .A2(new_n682), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n685));
  AOI211_X1 g260(.A(new_n681), .B(new_n683), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n684), .B2(new_n685), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT90), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT91), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1991), .B(G1996), .Z(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n689), .B(new_n690), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n696), .A2(new_n693), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n675), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n693), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n692), .A2(new_n694), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n699), .A2(new_n700), .A3(new_n674), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(G229));
  MUX2_X1   g277(.A(G24), .B(G290), .S(G16), .Z(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT92), .B(G1986), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n703), .A2(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(G29), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G25), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n475), .A2(G131), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n487), .A2(G119), .ZN(new_n711));
  OR2_X1    g286(.A1(G95), .A2(G2105), .ZN(new_n712));
  OAI211_X1 g287(.A(new_n712), .B(G2104), .C1(G107), .C2(new_n473), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n709), .B1(new_n715), .B2(new_n708), .ZN(new_n716));
  XOR2_X1   g291(.A(KEYINPUT35), .B(G1991), .Z(new_n717));
  XOR2_X1   g292(.A(new_n716), .B(new_n717), .Z(new_n718));
  NOR2_X1   g293(.A1(new_n707), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G16), .A2(G23), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT94), .Z(new_n721));
  INV_X1    g296(.A(G16), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(G288), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(KEYINPUT33), .B(G1976), .Z(new_n724));
  XNOR2_X1  g299(.A(new_n723), .B(new_n724), .ZN(new_n725));
  MUX2_X1   g300(.A(G6), .B(G305), .S(G16), .Z(new_n726));
  XOR2_X1   g301(.A(KEYINPUT32), .B(G1981), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n722), .A2(G22), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G166), .B2(new_n722), .ZN(new_n730));
  INV_X1    g305(.A(G1971), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n725), .A2(new_n728), .A3(new_n732), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT93), .B(KEYINPUT34), .Z(new_n734));
  OAI211_X1 g309(.A(new_n706), .B(new_n719), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(new_n734), .B2(new_n733), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT36), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n722), .A2(G20), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT23), .Z(new_n739));
  AOI21_X1  g314(.A(new_n739), .B1(G299), .B2(G16), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(G1956), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n708), .A2(G35), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G162), .B2(new_n708), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT29), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G2090), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT103), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n741), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(new_n746), .B2(new_n745), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT104), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n708), .A2(G26), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT28), .Z(new_n751));
  NAND2_X1  g326(.A1(new_n475), .A2(G140), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n487), .A2(G128), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n473), .A2(G116), .ZN(new_n754));
  OAI21_X1  g329(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n752), .B(new_n753), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n751), .B1(new_n756), .B2(G29), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT97), .B(G2067), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT31), .B(G11), .Z(new_n760));
  NOR2_X1   g335(.A1(new_n636), .A2(new_n708), .ZN(new_n761));
  INV_X1    g336(.A(G28), .ZN(new_n762));
  OR2_X1    g337(.A1(new_n762), .A2(KEYINPUT30), .ZN(new_n763));
  AOI21_X1  g338(.A(G29), .B1(new_n762), .B2(KEYINPUT30), .ZN(new_n764));
  AOI211_X1 g339(.A(new_n760), .B(new_n761), .C1(new_n763), .C2(new_n764), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n708), .A2(G32), .ZN(new_n766));
  NAND3_X1  g341(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT26), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n767), .A2(new_n768), .ZN(new_n770));
  AOI22_X1  g345(.A1(new_n769), .A2(new_n770), .B1(G105), .B2(new_n481), .ZN(new_n771));
  INV_X1    g346(.A(G141), .ZN(new_n772));
  INV_X1    g347(.A(G129), .ZN(new_n773));
  OAI221_X1 g348(.A(new_n771), .B1(new_n474), .B2(new_n772), .C1(new_n773), .C2(new_n486), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n766), .B1(new_n774), .B2(G29), .ZN(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT27), .B(G1996), .ZN(new_n776));
  OR2_X1    g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G34), .ZN(new_n778));
  AOI21_X1  g353(.A(G29), .B1(new_n778), .B2(KEYINPUT24), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(KEYINPUT24), .B2(new_n778), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n483), .B2(new_n708), .ZN(new_n781));
  INV_X1    g356(.A(G2084), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n781), .A2(new_n782), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n765), .A2(new_n777), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(G2072), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n708), .A2(G33), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT25), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n788), .B(new_n789), .ZN(new_n790));
  AOI22_X1  g365(.A1(new_n477), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n473), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(new_n475), .B2(G139), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n787), .B1(new_n793), .B2(new_n708), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT98), .Z(new_n795));
  AOI211_X1 g370(.A(new_n759), .B(new_n785), .C1(new_n786), .C2(new_n795), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n795), .A2(new_n786), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT99), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n722), .A2(G19), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n569), .B2(new_n722), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(G1341), .Z(new_n801));
  NAND3_X1  g376(.A1(new_n796), .A2(new_n798), .A3(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n744), .A2(G2090), .ZN(new_n803));
  INV_X1    g378(.A(G1961), .ZN(new_n804));
  NAND2_X1  g379(.A1(G171), .A2(G16), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G5), .B2(G16), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n775), .A2(new_n776), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT100), .ZN(new_n809));
  OAI211_X1 g384(.A(new_n807), .B(new_n809), .C1(new_n804), .C2(new_n806), .ZN(new_n810));
  NOR2_X1   g385(.A1(G16), .A2(G21), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n811), .B1(G168), .B2(G16), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(G1966), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n802), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  NOR2_X1   g389(.A1(G4), .A2(G16), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n815), .B1(new_n618), .B2(G16), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT95), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT96), .B(G1348), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n708), .A2(G27), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT101), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G164), .B2(new_n708), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT102), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G2078), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n749), .A2(new_n814), .A3(new_n819), .A4(new_n824), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n737), .A2(new_n825), .ZN(G311));
  XNOR2_X1  g401(.A(G311), .B(KEYINPUT105), .ZN(G150));
  NAND2_X1  g402(.A1(new_n618), .A2(G559), .ZN(new_n828));
  XOR2_X1   g403(.A(new_n828), .B(KEYINPUT38), .Z(new_n829));
  NAND2_X1  g404(.A1(new_n548), .A2(G67), .ZN(new_n830));
  INV_X1    g405(.A(G80), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(new_n525), .ZN(new_n832));
  AOI22_X1  g407(.A1(new_n832), .A2(G651), .B1(G55), .B2(new_n522), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT106), .B(G93), .Z(new_n834));
  NAND2_X1  g409(.A1(new_n556), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n568), .A2(new_n836), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n564), .A2(new_n833), .A3(new_n567), .A4(new_n835), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n829), .B(new_n840), .Z(new_n841));
  AND2_X1   g416(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n841), .A2(KEYINPUT39), .ZN(new_n843));
  NOR3_X1   g418(.A1(new_n842), .A2(new_n843), .A3(G860), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n836), .A2(G860), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n844), .A2(new_n846), .ZN(G145));
  XNOR2_X1  g422(.A(new_n636), .B(new_n483), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n491), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n793), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n756), .B(new_n774), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n640), .B(KEYINPUT107), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n475), .A2(G142), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n487), .A2(G130), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n473), .A2(G118), .ZN(new_n857));
  OAI21_X1  g432(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n858));
  OAI211_X1 g433(.A(new_n855), .B(new_n856), .C1(new_n857), .C2(new_n858), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT108), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n715), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n854), .B(new_n861), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n507), .A2(new_n497), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n862), .A2(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n862), .A2(new_n864), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n851), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n866), .A2(new_n851), .A3(new_n867), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n850), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(G37), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n866), .A2(new_n867), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(new_n793), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n874), .A2(new_n849), .A3(new_n868), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n871), .A2(new_n872), .A3(new_n875), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g452(.A(KEYINPUT112), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n840), .B(new_n628), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n611), .A2(new_n613), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n617), .A2(new_n616), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(G299), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n618), .A2(G299), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n879), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(KEYINPUT109), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(KEYINPUT110), .A3(new_n883), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT110), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n889), .B1(new_n618), .B2(G299), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n888), .A2(new_n890), .A3(new_n885), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n884), .A2(new_n885), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT111), .B1(new_n894), .B2(new_n892), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT111), .ZN(new_n896));
  NAND4_X1  g471(.A1(new_n884), .A2(new_n885), .A3(new_n896), .A4(KEYINPUT41), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n879), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n878), .B1(new_n887), .B2(new_n899), .ZN(new_n900));
  XOR2_X1   g475(.A(G288), .B(G305), .Z(new_n901));
  XNOR2_X1  g476(.A(G290), .B(G166), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n901), .B(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n903), .B(KEYINPUT42), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n887), .A2(new_n878), .A3(new_n899), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n900), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  AOI211_X1 g482(.A(new_n878), .B(new_n904), .C1(new_n887), .C2(new_n899), .ZN(new_n908));
  OAI21_X1  g483(.A(G868), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n836), .A2(new_n622), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(G295));
  NAND2_X1  g486(.A1(new_n909), .A2(new_n910), .ZN(G331));
  INV_X1    g487(.A(KEYINPUT44), .ZN(new_n913));
  OAI21_X1  g488(.A(G286), .B1(new_n837), .B2(new_n839), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n568), .A2(new_n836), .ZN(new_n915));
  NAND3_X1  g490(.A1(G168), .A2(new_n915), .A3(new_n838), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(G301), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(G171), .A3(new_n916), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n918), .A2(new_n894), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT113), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n919), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n921), .B1(new_n898), .B2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT113), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n898), .A2(new_n924), .A3(new_n922), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n903), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n898), .A2(new_n922), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(KEYINPUT113), .A3(new_n920), .ZN(new_n930));
  INV_X1    g505(.A(new_n903), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n930), .A2(new_n931), .A3(new_n925), .ZN(new_n932));
  NAND4_X1  g507(.A1(new_n927), .A2(new_n928), .A3(new_n872), .A4(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n892), .B1(new_n918), .B2(new_n919), .ZN(new_n934));
  OR2_X1    g509(.A1(new_n934), .A2(new_n894), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n903), .B1(new_n934), .B2(new_n891), .ZN(new_n936));
  AOI21_X1  g511(.A(G37), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n931), .B1(new_n930), .B2(new_n925), .ZN(new_n939));
  OAI21_X1  g514(.A(KEYINPUT43), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n913), .B1(new_n933), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n927), .A2(new_n872), .A3(new_n932), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n942), .A2(KEYINPUT43), .B1(new_n943), .B2(new_n937), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n941), .B1(new_n944), .B2(new_n913), .ZN(G397));
  INV_X1    g520(.A(KEYINPUT124), .ZN(new_n946));
  INV_X1    g521(.A(G8), .ZN(new_n947));
  INV_X1    g522(.A(new_n497), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n465), .A2(KEYINPUT67), .A3(new_n463), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT67), .B1(new_n469), .B2(G2104), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n469), .A2(KEYINPUT66), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n950), .B1(new_n953), .B2(G2104), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n503), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n955), .A2(new_n505), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n472), .A2(KEYINPUT68), .A3(new_n503), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT69), .B1(new_n958), .B2(new_n501), .ZN(new_n959));
  INV_X1    g534(.A(new_n510), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n948), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT118), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(G1384), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n964), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT118), .B1(G164), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n476), .A2(G40), .A3(new_n482), .ZN(new_n968));
  INV_X1    g543(.A(G1384), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n507), .B2(new_n497), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n968), .B1(new_n970), .B2(new_n963), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n965), .A2(new_n967), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1966), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n975));
  INV_X1    g550(.A(new_n968), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n976), .B1(new_n970), .B2(KEYINPUT50), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n978), .A3(new_n782), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n947), .B1(new_n974), .B2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT116), .B(G8), .ZN(new_n981));
  NOR2_X1   g556(.A1(G168), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT51), .B1(new_n980), .B2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n982), .A2(KEYINPUT51), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n961), .A2(new_n969), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n977), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n973), .A2(new_n972), .B1(new_n986), .B2(new_n782), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n984), .B1(new_n987), .B2(new_n981), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n983), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n982), .ZN(new_n990));
  NOR2_X1   g565(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n946), .B1(new_n989), .B2(new_n992), .ZN(new_n993));
  AOI211_X1 g568(.A(KEYINPUT124), .B(new_n991), .C1(new_n983), .C2(new_n988), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT62), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n990), .B1(new_n987), .B2(new_n947), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n974), .A2(new_n979), .ZN(new_n997));
  INV_X1    g572(.A(new_n981), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  AOI22_X1  g574(.A1(new_n996), .A2(KEYINPUT51), .B1(new_n999), .B2(new_n984), .ZN(new_n1000));
  OAI21_X1  g575(.A(KEYINPUT124), .B1(new_n1000), .B2(new_n991), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT62), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n989), .A2(new_n946), .A3(new_n992), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  XOR2_X1   g579(.A(KEYINPUT117), .B(G86), .Z(new_n1005));
  NAND2_X1  g580(.A1(new_n556), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n593), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(G1981), .ZN(new_n1008));
  OR2_X1    g583(.A1(G305), .A2(G1981), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1008), .A2(KEYINPUT49), .A3(new_n1009), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n500), .B1(new_n956), .B2(new_n957), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1384), .B1(new_n1011), .B2(new_n948), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n981), .B1(new_n1012), .B2(new_n976), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT49), .ZN(new_n1014));
  INV_X1    g589(.A(G1981), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1015), .B1(new_n1006), .B2(new_n593), .ZN(new_n1016));
  NOR2_X1   g591(.A1(G305), .A2(G1981), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n1014), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1010), .A2(new_n1013), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(G288), .B2(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n588), .A2(new_n587), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1022), .A2(G1976), .A3(new_n584), .A4(new_n585), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1021), .A2(new_n1013), .A3(new_n1023), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1013), .B1(G288), .B2(new_n1020), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(KEYINPUT52), .ZN(new_n1026));
  AND3_X1   g601(.A1(new_n1019), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G303), .A2(G8), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT55), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT115), .B(G2090), .Z(new_n1031));
  AND3_X1   g606(.A1(new_n975), .A2(new_n978), .A3(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n963), .B1(G164), .B2(G1384), .ZN(new_n1033));
  XNOR2_X1  g608(.A(KEYINPUT114), .B(G1384), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n863), .A2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n968), .B1(new_n1035), .B2(KEYINPUT45), .ZN(new_n1036));
  AOI21_X1  g611(.A(G1971), .B1(new_n1033), .B2(new_n1036), .ZN(new_n1037));
  OAI211_X1 g612(.A(new_n1030), .B(G8), .C1(new_n1032), .C2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT50), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n976), .B1(new_n1012), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G164), .A2(G1384), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1041), .B2(new_n1039), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1042), .A2(new_n1031), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1033), .A2(new_n1036), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1044), .A2(new_n731), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n981), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1027), .B(new_n1038), .C1(new_n1030), .C2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  INV_X1    g624(.A(G2078), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n965), .A2(new_n967), .A3(new_n1050), .A4(new_n971), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT125), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1049), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n1052), .B2(new_n1051), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1033), .A2(new_n1036), .A3(new_n1050), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n975), .A2(new_n978), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1055), .A2(new_n1049), .B1(new_n1056), .B2(new_n804), .ZN(new_n1057));
  AOI21_X1  g632(.A(G301), .B1(new_n1054), .B2(new_n1057), .ZN(new_n1058));
  AND2_X1   g633(.A1(new_n1048), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n995), .A2(new_n1004), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT127), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT127), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n995), .A2(new_n1004), .A3(new_n1062), .A4(new_n1059), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n997), .A2(G168), .A3(new_n998), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1064), .B1(new_n1047), .B2(new_n1065), .ZN(new_n1066));
  OAI21_X1  g641(.A(G8), .B1(new_n1032), .B2(new_n1037), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1064), .B1(new_n1067), .B2(new_n1029), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1068), .A2(new_n1038), .A3(new_n1027), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1066), .B1(new_n1065), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1038), .ZN(new_n1071));
  NOR2_X1   g646(.A1(G288), .A2(G1976), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1019), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(new_n1009), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1071), .A2(new_n1027), .B1(new_n1074), .B2(new_n1013), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1070), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT57), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1077), .A2(KEYINPUT57), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(G299), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  AND2_X1   g656(.A1(new_n578), .A2(new_n580), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1082), .A2(KEYINPUT119), .A3(new_n1083), .A4(new_n577), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1081), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1042), .A2(G1956), .ZN(new_n1086));
  XNOR2_X1  g661(.A(KEYINPUT56), .B(G2072), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1033), .A2(new_n1036), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1085), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1085), .ZN(new_n1091));
  OAI211_X1 g666(.A(new_n1091), .B(new_n1088), .C1(new_n1042), .C2(G1956), .ZN(new_n1092));
  AOI21_X1  g667(.A(KEYINPUT61), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT60), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1012), .A2(new_n976), .ZN(new_n1095));
  INV_X1    g670(.A(new_n818), .ZN(new_n1096));
  OAI221_X1 g671(.A(new_n882), .B1(G2067), .B2(new_n1095), .C1(new_n986), .C2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(new_n1096), .B1(new_n975), .B2(new_n978), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1095), .A2(G2067), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n618), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1094), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  NOR4_X1   g676(.A1(new_n1098), .A2(new_n882), .A3(KEYINPUT60), .A4(new_n1099), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1093), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT122), .B1(new_n1044), .B2(G1996), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n1105));
  INV_X1    g680(.A(G1996), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1033), .A2(new_n1036), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT58), .B(G1341), .Z(new_n1108));
  NAND2_X1  g683(.A1(new_n1095), .A2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1104), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(new_n569), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT59), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(new_n1113), .A3(new_n569), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT123), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1092), .A2(KEYINPUT61), .ZN(new_n1117));
  INV_X1    g692(.A(G1956), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n985), .A2(KEYINPUT50), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1118), .B1(new_n1119), .B2(new_n1040), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1085), .A2(KEYINPUT120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1081), .A2(new_n1084), .A3(new_n1122), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1120), .A2(new_n1088), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1116), .B1(new_n1117), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1086), .B2(new_n1089), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1127), .A2(KEYINPUT123), .A3(KEYINPUT61), .A4(new_n1092), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1125), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1103), .A2(new_n1115), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1100), .ZN(new_n1131));
  OAI211_X1 g706(.A(KEYINPUT121), .B(new_n1092), .C1(new_n1124), .C2(new_n1131), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1127), .A2(new_n1100), .ZN(new_n1134));
  AOI21_X1  g709(.A(KEYINPUT121), .B1(new_n1134), .B2(new_n1092), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1130), .A2(new_n1136), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1054), .A2(G301), .A3(new_n1057), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(KEYINPUT126), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT126), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n1054), .A2(new_n1140), .A3(G301), .A4(new_n1057), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n963), .B1(new_n863), .B2(new_n1034), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1036), .A2(KEYINPUT53), .A3(new_n1050), .A4(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1057), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1142), .B1(new_n1145), .B2(G171), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1139), .A2(new_n1141), .A3(new_n1146), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1145), .A2(G171), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1142), .B1(new_n1058), .B2(new_n1148), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1147), .A2(new_n1048), .A3(new_n1149), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1076), .B1(new_n1137), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1061), .A2(new_n1063), .A3(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1143), .A2(new_n968), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n756), .B(G2067), .Z(new_n1154));
  XNOR2_X1  g729(.A(new_n774), .B(new_n1106), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  XOR2_X1   g731(.A(new_n714), .B(new_n717), .Z(new_n1157));
  NOR2_X1   g732(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(G290), .B(G1986), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1153), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1152), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1154), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1153), .B1(new_n1163), .B2(new_n774), .ZN(new_n1164));
  NOR4_X1   g739(.A1(new_n1143), .A2(KEYINPUT46), .A3(G1996), .A4(new_n968), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT46), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1166), .B1(new_n1153), .B2(new_n1106), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n1164), .B1(new_n1165), .B2(new_n1167), .ZN(new_n1168));
  XNOR2_X1  g743(.A(new_n1168), .B(KEYINPUT47), .ZN(new_n1169));
  NOR2_X1   g744(.A1(G290), .A2(G1986), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1153), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1159), .A2(new_n1153), .B1(new_n1172), .B2(KEYINPUT48), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n1173), .B1(KEYINPUT48), .B2(new_n1172), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n715), .A2(new_n717), .ZN(new_n1175));
  OAI22_X1  g750(.A1(new_n1156), .A2(new_n1175), .B1(G2067), .B2(new_n756), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(new_n1153), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1169), .A2(new_n1174), .A3(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1162), .A2(new_n1178), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g754(.A1(new_n660), .A2(new_n460), .A3(G227), .ZN(new_n1181));
  INV_X1    g755(.A(new_n1181), .ZN(new_n1182));
  AND3_X1   g756(.A1(new_n698), .A2(new_n701), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g757(.A1(new_n1183), .A2(new_n876), .ZN(new_n1184));
  NOR2_X1   g758(.A1(new_n1184), .A2(new_n944), .ZN(G308));
  AND2_X1   g759(.A1(new_n942), .A2(KEYINPUT43), .ZN(new_n1186));
  NOR3_X1   g760(.A1(new_n938), .A2(new_n939), .A3(KEYINPUT43), .ZN(new_n1187));
  OAI211_X1 g761(.A(new_n876), .B(new_n1183), .C1(new_n1186), .C2(new_n1187), .ZN(G225));
endmodule


