

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584;

  INV_X1 U320 ( .A(KEYINPUT69), .ZN(n430) );
  XNOR2_X1 U321 ( .A(n418), .B(KEYINPUT104), .ZN(n419) );
  XOR2_X1 U322 ( .A(KEYINPUT93), .B(n376), .Z(n548) );
  XOR2_X1 U323 ( .A(n301), .B(n300), .Z(n288) );
  XOR2_X1 U324 ( .A(n573), .B(KEYINPUT59), .Z(n289) );
  INV_X1 U325 ( .A(KEYINPUT46), .ZN(n504) );
  NOR2_X1 U326 ( .A1(n538), .A2(n508), .ZN(n509) );
  XNOR2_X1 U327 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U328 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U329 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U330 ( .A(n429), .B(n428), .ZN(n436) );
  XNOR2_X1 U331 ( .A(n302), .B(n288), .ZN(n303) );
  XNOR2_X1 U332 ( .A(n436), .B(n435), .ZN(n438) );
  XNOR2_X1 U333 ( .A(n420), .B(n419), .ZN(n493) );
  XNOR2_X1 U334 ( .A(n304), .B(n303), .ZN(n305) );
  NOR2_X1 U335 ( .A1(n569), .A2(n568), .ZN(n581) );
  INV_X1 U336 ( .A(G43GAT), .ZN(n458) );
  XNOR2_X1 U337 ( .A(n458), .B(KEYINPUT40), .ZN(n459) );
  XNOR2_X1 U338 ( .A(n460), .B(n459), .ZN(G1330GAT) );
  NAND2_X1 U339 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XOR2_X1 U340 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n291) );
  XNOR2_X1 U341 ( .A(G43GAT), .B(G190GAT), .ZN(n290) );
  XNOR2_X1 U342 ( .A(n291), .B(n290), .ZN(n293) );
  XOR2_X1 U343 ( .A(G99GAT), .B(G134GAT), .Z(n292) );
  XNOR2_X1 U344 ( .A(n293), .B(n292), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n306) );
  XOR2_X1 U346 ( .A(KEYINPUT84), .B(KEYINPUT17), .Z(n297) );
  XNOR2_X1 U347 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n298) );
  XNOR2_X1 U349 ( .A(KEYINPUT19), .B(n298), .ZN(n346) );
  XOR2_X1 U350 ( .A(G169GAT), .B(n346), .Z(n304) );
  XNOR2_X1 U351 ( .A(G127GAT), .B(KEYINPUT82), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n299), .B(KEYINPUT0), .ZN(n326) );
  XOR2_X1 U353 ( .A(G176GAT), .B(n326), .Z(n302) );
  XOR2_X1 U354 ( .A(G120GAT), .B(G71GAT), .Z(n301) );
  XNOR2_X1 U355 ( .A(G15GAT), .B(G113GAT), .ZN(n300) );
  XNOR2_X1 U356 ( .A(n306), .B(n305), .ZN(n552) );
  XOR2_X1 U357 ( .A(KEYINPUT90), .B(KEYINPUT5), .Z(n308) );
  XOR2_X1 U358 ( .A(G113GAT), .B(G1GAT), .Z(n422) );
  XOR2_X1 U359 ( .A(G134GAT), .B(G162GAT), .Z(n407) );
  XNOR2_X1 U360 ( .A(n422), .B(n407), .ZN(n307) );
  XOR2_X1 U361 ( .A(n308), .B(n307), .Z(n318) );
  INV_X1 U362 ( .A(KEYINPUT2), .ZN(n309) );
  NAND2_X1 U363 ( .A1(G155GAT), .A2(n309), .ZN(n312) );
  INV_X1 U364 ( .A(G155GAT), .ZN(n310) );
  NAND2_X1 U365 ( .A1(n310), .A2(KEYINPUT2), .ZN(n311) );
  NAND2_X1 U366 ( .A1(n312), .A2(n311), .ZN(n314) );
  XNOR2_X1 U367 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n354) );
  XOR2_X1 U369 ( .A(n354), .B(KEYINPUT91), .Z(n316) );
  NAND2_X1 U370 ( .A1(G225GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U371 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U372 ( .A(n318), .B(n317), .ZN(n320) );
  XNOR2_X1 U373 ( .A(G29GAT), .B(G85GAT), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n320), .B(n319), .ZN(n324) );
  XOR2_X1 U375 ( .A(KEYINPUT4), .B(KEYINPUT92), .Z(n322) );
  XNOR2_X1 U376 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n321) );
  XNOR2_X1 U377 ( .A(n322), .B(n321), .ZN(n323) );
  XOR2_X1 U378 ( .A(n324), .B(n323), .Z(n328) );
  XNOR2_X1 U379 ( .A(G120GAT), .B(G148GAT), .ZN(n325) );
  XNOR2_X1 U380 ( .A(n325), .B(G57GAT), .ZN(n448) );
  XNOR2_X1 U381 ( .A(n326), .B(n448), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n376) );
  XOR2_X1 U383 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n330) );
  XNOR2_X1 U384 ( .A(KEYINPUT88), .B(KEYINPUT21), .ZN(n329) );
  XNOR2_X1 U385 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U386 ( .A(n331), .B(G211GAT), .Z(n333) );
  XNOR2_X1 U387 ( .A(G197GAT), .B(G204GAT), .ZN(n332) );
  XNOR2_X1 U388 ( .A(n333), .B(n332), .ZN(n362) );
  INV_X1 U389 ( .A(G218GAT), .ZN(n334) );
  NAND2_X1 U390 ( .A1(G92GAT), .A2(n334), .ZN(n337) );
  INV_X1 U391 ( .A(G92GAT), .ZN(n335) );
  NAND2_X1 U392 ( .A1(n335), .A2(G218GAT), .ZN(n336) );
  NAND2_X1 U393 ( .A1(n337), .A2(n336), .ZN(n339) );
  XNOR2_X1 U394 ( .A(G36GAT), .B(G190GAT), .ZN(n338) );
  XNOR2_X1 U395 ( .A(n339), .B(n338), .ZN(n408) );
  XOR2_X1 U396 ( .A(G176GAT), .B(G64GAT), .Z(n450) );
  XNOR2_X1 U397 ( .A(n408), .B(n450), .ZN(n341) );
  AND2_X1 U398 ( .A1(G226GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U400 ( .A(n342), .B(KEYINPUT95), .ZN(n344) );
  XOR2_X1 U401 ( .A(G169GAT), .B(G8GAT), .Z(n421) );
  XOR2_X1 U402 ( .A(n421), .B(KEYINPUT94), .Z(n343) );
  XNOR2_X1 U403 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U404 ( .A(n362), .B(n345), .Z(n347) );
  XNOR2_X1 U405 ( .A(n347), .B(n346), .ZN(n542) );
  XOR2_X1 U406 ( .A(KEYINPUT27), .B(KEYINPUT96), .Z(n348) );
  XOR2_X1 U407 ( .A(n542), .B(n348), .Z(n368) );
  NOR2_X1 U408 ( .A1(n548), .A2(n368), .ZN(n517) );
  NAND2_X1 U409 ( .A1(n552), .A2(n517), .ZN(n365) );
  XOR2_X1 U410 ( .A(G148GAT), .B(G106GAT), .Z(n350) );
  XNOR2_X1 U411 ( .A(G22GAT), .B(G218GAT), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U413 ( .A(n351), .B(G162GAT), .Z(n353) );
  XOR2_X1 U414 ( .A(KEYINPUT74), .B(G78GAT), .Z(n451) );
  XNOR2_X1 U415 ( .A(G50GAT), .B(n451), .ZN(n352) );
  XNOR2_X1 U416 ( .A(n353), .B(n352), .ZN(n358) );
  XOR2_X1 U417 ( .A(KEYINPUT22), .B(n354), .Z(n356) );
  NAND2_X1 U418 ( .A1(G228GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U419 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U420 ( .A(n358), .B(n357), .Z(n364) );
  XOR2_X1 U421 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n360) );
  XNOR2_X1 U422 ( .A(KEYINPUT85), .B(KEYINPUT89), .ZN(n359) );
  XNOR2_X1 U423 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U425 ( .A(n364), .B(n363), .ZN(n549) );
  XNOR2_X1 U426 ( .A(n549), .B(KEYINPUT28), .ZN(n520) );
  NOR2_X1 U427 ( .A1(n365), .A2(n520), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n366), .B(KEYINPUT97), .ZN(n378) );
  NAND2_X1 U429 ( .A1(n552), .A2(n549), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n367), .B(KEYINPUT26), .ZN(n569) );
  NOR2_X1 U431 ( .A1(n569), .A2(n368), .ZN(n370) );
  INV_X1 U432 ( .A(KEYINPUT98), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n370), .B(n369), .ZN(n374) );
  NOR2_X1 U434 ( .A1(n552), .A2(n542), .ZN(n371) );
  NOR2_X1 U435 ( .A1(n549), .A2(n371), .ZN(n372) );
  XNOR2_X1 U436 ( .A(KEYINPUT25), .B(n372), .ZN(n373) );
  NAND2_X1 U437 ( .A1(n374), .A2(n373), .ZN(n375) );
  NAND2_X1 U438 ( .A1(n376), .A2(n375), .ZN(n377) );
  NAND2_X1 U439 ( .A1(n378), .A2(n377), .ZN(n379) );
  XNOR2_X1 U440 ( .A(KEYINPUT99), .B(n379), .ZN(n464) );
  XOR2_X1 U441 ( .A(KEYINPUT14), .B(KEYINPUT78), .Z(n381) );
  XNOR2_X1 U442 ( .A(G1GAT), .B(KEYINPUT15), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n399) );
  XOR2_X1 U444 ( .A(KEYINPUT79), .B(G78GAT), .Z(n383) );
  XNOR2_X1 U445 ( .A(G183GAT), .B(G127GAT), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U447 ( .A(KEYINPUT80), .B(G57GAT), .Z(n385) );
  XNOR2_X1 U448 ( .A(G8GAT), .B(G64GAT), .ZN(n384) );
  XNOR2_X1 U449 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U450 ( .A(n387), .B(n386), .Z(n393) );
  XNOR2_X1 U451 ( .A(G22GAT), .B(G15GAT), .ZN(n388) );
  XNOR2_X1 U452 ( .A(n388), .B(KEYINPUT68), .ZN(n433) );
  XOR2_X1 U453 ( .A(G155GAT), .B(G211GAT), .Z(n390) );
  NAND2_X1 U454 ( .A1(G231GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U455 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U456 ( .A(n433), .B(n391), .ZN(n392) );
  XNOR2_X1 U457 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U458 ( .A(n394), .B(KEYINPUT81), .Z(n397) );
  XNOR2_X1 U459 ( .A(G71GAT), .B(KEYINPUT71), .ZN(n395) );
  XNOR2_X1 U460 ( .A(n395), .B(KEYINPUT13), .ZN(n444) );
  XNOR2_X1 U461 ( .A(n444), .B(KEYINPUT12), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U463 ( .A(n399), .B(n398), .ZN(n579) );
  NOR2_X1 U464 ( .A1(n464), .A2(n579), .ZN(n400) );
  XNOR2_X1 U465 ( .A(KEYINPUT102), .B(n400), .ZN(n417) );
  XOR2_X1 U466 ( .A(KEYINPUT8), .B(G50GAT), .Z(n402) );
  XNOR2_X1 U467 ( .A(G43GAT), .B(G29GAT), .ZN(n401) );
  XNOR2_X1 U468 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U469 ( .A(KEYINPUT7), .B(n403), .ZN(n437) );
  XOR2_X1 U470 ( .A(KEYINPUT11), .B(KEYINPUT75), .Z(n405) );
  XNOR2_X1 U471 ( .A(KEYINPUT64), .B(KEYINPUT10), .ZN(n404) );
  XNOR2_X1 U472 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U473 ( .A(n437), .B(n406), .Z(n416) );
  XOR2_X1 U474 ( .A(n408), .B(n407), .Z(n410) );
  NAND2_X1 U475 ( .A1(G232GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U476 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U477 ( .A(n411), .B(KEYINPUT9), .Z(n414) );
  XNOR2_X1 U478 ( .A(G99GAT), .B(G106GAT), .ZN(n412) );
  XNOR2_X1 U479 ( .A(n412), .B(G85GAT), .ZN(n445) );
  XNOR2_X1 U480 ( .A(n445), .B(KEYINPUT76), .ZN(n413) );
  XNOR2_X1 U481 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U482 ( .A(n416), .B(n415), .ZN(n538) );
  XOR2_X1 U483 ( .A(KEYINPUT77), .B(n538), .Z(n564) );
  XNOR2_X1 U484 ( .A(KEYINPUT36), .B(n564), .ZN(n582) );
  NAND2_X1 U485 ( .A1(n417), .A2(n582), .ZN(n420) );
  XOR2_X1 U486 ( .A(KEYINPUT37), .B(KEYINPUT103), .Z(n418) );
  XOR2_X1 U487 ( .A(KEYINPUT29), .B(G141GAT), .Z(n424) );
  XNOR2_X1 U488 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U489 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U490 ( .A(n425), .B(G197GAT), .Z(n429) );
  XOR2_X1 U491 ( .A(KEYINPUT65), .B(KEYINPUT67), .Z(n427) );
  XNOR2_X1 U492 ( .A(KEYINPUT66), .B(KEYINPUT30), .ZN(n426) );
  XNOR2_X1 U493 ( .A(n427), .B(n426), .ZN(n428) );
  NAND2_X1 U494 ( .A1(G229GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n434), .B(G36GAT), .ZN(n435) );
  XOR2_X1 U496 ( .A(n438), .B(n437), .Z(n570) );
  XNOR2_X1 U497 ( .A(n570), .B(KEYINPUT70), .ZN(n553) );
  INV_X1 U498 ( .A(n553), .ZN(n456) );
  XOR2_X1 U499 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n440) );
  XNOR2_X1 U500 ( .A(G204GAT), .B(G92GAT), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n455) );
  XOR2_X1 U502 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n442) );
  NAND2_X1 U503 ( .A1(G230GAT), .A2(G233GAT), .ZN(n441) );
  XNOR2_X1 U504 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U505 ( .A(n443), .B(KEYINPUT31), .Z(n447) );
  XNOR2_X1 U506 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U507 ( .A(n447), .B(n446), .ZN(n449) );
  XOR2_X1 U508 ( .A(n449), .B(n448), .Z(n453) );
  XNOR2_X1 U509 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U510 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U511 ( .A(n455), .B(n454), .ZN(n575) );
  NOR2_X1 U512 ( .A1(n456), .A2(n575), .ZN(n465) );
  NAND2_X1 U513 ( .A1(n493), .A2(n465), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n457), .B(KEYINPUT38), .ZN(n478) );
  NOR2_X1 U515 ( .A1(n552), .A2(n478), .ZN(n460) );
  INV_X1 U516 ( .A(n579), .ZN(n461) );
  NOR2_X1 U517 ( .A1(n564), .A2(n461), .ZN(n462) );
  XOR2_X1 U518 ( .A(KEYINPUT16), .B(n462), .Z(n463) );
  NOR2_X1 U519 ( .A1(n464), .A2(n463), .ZN(n482) );
  NAND2_X1 U520 ( .A1(n465), .A2(n482), .ZN(n472) );
  NOR2_X1 U521 ( .A1(n548), .A2(n472), .ZN(n466) );
  XOR2_X1 U522 ( .A(KEYINPUT34), .B(n466), .Z(n467) );
  XNOR2_X1 U523 ( .A(G1GAT), .B(n467), .ZN(G1324GAT) );
  NOR2_X1 U524 ( .A1(n542), .A2(n472), .ZN(n468) );
  XOR2_X1 U525 ( .A(G8GAT), .B(n468), .Z(G1325GAT) );
  NOR2_X1 U526 ( .A1(n552), .A2(n472), .ZN(n470) );
  XNOR2_X1 U527 ( .A(KEYINPUT35), .B(KEYINPUT100), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U529 ( .A(G15GAT), .B(n471), .ZN(G1326GAT) );
  INV_X1 U530 ( .A(n520), .ZN(n499) );
  NOR2_X1 U531 ( .A1(n499), .A2(n472), .ZN(n474) );
  XNOR2_X1 U532 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n474), .B(n473), .ZN(G1327GAT) );
  XNOR2_X1 U534 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n476) );
  NOR2_X1 U535 ( .A1(n548), .A2(n478), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n476), .B(n475), .ZN(G1328GAT) );
  NOR2_X1 U537 ( .A1(n542), .A2(n478), .ZN(n477) );
  XOR2_X1 U538 ( .A(G36GAT), .B(n477), .Z(G1329GAT) );
  NOR2_X1 U539 ( .A1(n499), .A2(n478), .ZN(n479) );
  XOR2_X1 U540 ( .A(G50GAT), .B(n479), .Z(G1331GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n481) );
  XNOR2_X1 U542 ( .A(G57GAT), .B(KEYINPUT105), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(n484) );
  XNOR2_X1 U544 ( .A(KEYINPUT41), .B(n575), .ZN(n503) );
  NOR2_X1 U545 ( .A1(n570), .A2(n503), .ZN(n494) );
  NAND2_X1 U546 ( .A1(n494), .A2(n482), .ZN(n488) );
  NOR2_X1 U547 ( .A1(n548), .A2(n488), .ZN(n483) );
  XOR2_X1 U548 ( .A(n484), .B(n483), .Z(G1332GAT) );
  NOR2_X1 U549 ( .A1(n542), .A2(n488), .ZN(n486) );
  XNOR2_X1 U550 ( .A(G64GAT), .B(KEYINPUT107), .ZN(n485) );
  XNOR2_X1 U551 ( .A(n486), .B(n485), .ZN(G1333GAT) );
  NOR2_X1 U552 ( .A1(n552), .A2(n488), .ZN(n487) );
  XOR2_X1 U553 ( .A(G71GAT), .B(n487), .Z(G1334GAT) );
  NOR2_X1 U554 ( .A1(n488), .A2(n499), .ZN(n492) );
  XOR2_X1 U555 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n490) );
  XNOR2_X1 U556 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n489) );
  XNOR2_X1 U557 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U558 ( .A(n492), .B(n491), .ZN(G1335GAT) );
  NAND2_X1 U559 ( .A1(n494), .A2(n493), .ZN(n498) );
  NOR2_X1 U560 ( .A1(n548), .A2(n498), .ZN(n495) );
  XOR2_X1 U561 ( .A(G85GAT), .B(n495), .Z(G1336GAT) );
  NOR2_X1 U562 ( .A1(n542), .A2(n498), .ZN(n496) );
  XOR2_X1 U563 ( .A(G92GAT), .B(n496), .Z(G1337GAT) );
  NOR2_X1 U564 ( .A1(n552), .A2(n498), .ZN(n497) );
  XOR2_X1 U565 ( .A(G99GAT), .B(n497), .Z(G1338GAT) );
  NOR2_X1 U566 ( .A1(n499), .A2(n498), .ZN(n501) );
  XNOR2_X1 U567 ( .A(KEYINPUT110), .B(KEYINPUT44), .ZN(n500) );
  XNOR2_X1 U568 ( .A(n501), .B(n500), .ZN(n502) );
  XOR2_X1 U569 ( .A(G106GAT), .B(n502), .Z(G1339GAT) );
  INV_X1 U570 ( .A(n503), .ZN(n559) );
  NAND2_X1 U571 ( .A1(n559), .A2(n570), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n505), .B(n504), .ZN(n506) );
  NOR2_X1 U573 ( .A1(n579), .A2(n506), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n507), .B(KEYINPUT111), .ZN(n508) );
  XNOR2_X1 U575 ( .A(KEYINPUT47), .B(n509), .ZN(n515) );
  XOR2_X1 U576 ( .A(KEYINPUT45), .B(KEYINPUT112), .Z(n511) );
  NAND2_X1 U577 ( .A1(n579), .A2(n582), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n511), .B(n510), .ZN(n513) );
  NOR2_X1 U579 ( .A1(n553), .A2(n575), .ZN(n512) );
  NAND2_X1 U580 ( .A1(n513), .A2(n512), .ZN(n514) );
  NAND2_X1 U581 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(KEYINPUT48), .B(n516), .ZN(n544) );
  NAND2_X1 U583 ( .A1(n544), .A2(n517), .ZN(n531) );
  NOR2_X1 U584 ( .A1(n552), .A2(n531), .ZN(n518) );
  XNOR2_X1 U585 ( .A(n518), .B(KEYINPUT113), .ZN(n519) );
  NOR2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n527) );
  NAND2_X1 U587 ( .A1(n527), .A2(n553), .ZN(n521) );
  XNOR2_X1 U588 ( .A(G113GAT), .B(n521), .ZN(G1340GAT) );
  XOR2_X1 U589 ( .A(G120GAT), .B(KEYINPUT49), .Z(n523) );
  NAND2_X1 U590 ( .A1(n527), .A2(n559), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(G1341GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n525) );
  NAND2_X1 U593 ( .A1(n527), .A2(n579), .ZN(n524) );
  XNOR2_X1 U594 ( .A(n525), .B(n524), .ZN(n526) );
  XOR2_X1 U595 ( .A(G127GAT), .B(n526), .Z(G1342GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT51), .B(KEYINPUT115), .Z(n529) );
  NAND2_X1 U597 ( .A1(n527), .A2(n564), .ZN(n528) );
  XNOR2_X1 U598 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U599 ( .A(G134GAT), .B(n530), .Z(G1343GAT) );
  XNOR2_X1 U600 ( .A(G141GAT), .B(KEYINPUT116), .ZN(n533) );
  NOR2_X1 U601 ( .A1(n569), .A2(n531), .ZN(n539) );
  NAND2_X1 U602 ( .A1(n570), .A2(n539), .ZN(n532) );
  XNOR2_X1 U603 ( .A(n533), .B(n532), .ZN(G1344GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n535) );
  NAND2_X1 U605 ( .A1(n539), .A2(n559), .ZN(n534) );
  XNOR2_X1 U606 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U607 ( .A(G148GAT), .B(n536), .ZN(G1345GAT) );
  NAND2_X1 U608 ( .A1(n579), .A2(n539), .ZN(n537) );
  XNOR2_X1 U609 ( .A(n537), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U610 ( .A(G162GAT), .B(KEYINPUT117), .Z(n541) );
  NAND2_X1 U611 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U612 ( .A(n541), .B(n540), .ZN(G1347GAT) );
  XOR2_X1 U613 ( .A(KEYINPUT118), .B(n542), .Z(n543) );
  NAND2_X1 U614 ( .A1(n544), .A2(n543), .ZN(n546) );
  XNOR2_X1 U615 ( .A(KEYINPUT119), .B(KEYINPUT54), .ZN(n545) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n568) );
  NOR2_X1 U617 ( .A1(n549), .A2(n568), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n550), .B(KEYINPUT55), .ZN(n551) );
  NOR2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n565) );
  NAND2_X1 U620 ( .A1(n553), .A2(n565), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n554), .B(KEYINPUT120), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G169GAT), .B(n555), .ZN(G1348GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n557) );
  XNOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n556) );
  XNOR2_X1 U625 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U626 ( .A(KEYINPUT121), .B(n558), .Z(n561) );
  NAND2_X1 U627 ( .A1(n565), .A2(n559), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  XOR2_X1 U629 ( .A(G183GAT), .B(KEYINPUT123), .Z(n563) );
  NAND2_X1 U630 ( .A1(n565), .A2(n579), .ZN(n562) );
  XNOR2_X1 U631 ( .A(n563), .B(n562), .ZN(G1350GAT) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(KEYINPUT58), .ZN(n567) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(n567), .ZN(G1351GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n572) );
  NAND2_X1 U636 ( .A1(n581), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n574) );
  XNOR2_X1 U639 ( .A(n289), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U640 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n577) );
  NAND2_X1 U641 ( .A1(n581), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G204GAT), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n581), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

