//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n762, new_n763, new_n764,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070;
  XNOR2_X1  g000(.A(KEYINPUT70), .B(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G140), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G125), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n192), .A2(G140), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT16), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n194), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n194), .A2(new_n197), .A3(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT23), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G128), .ZN(new_n205));
  INV_X1    g019(.A(G128), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT23), .A3(G119), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n205), .B(new_n207), .C1(G119), .C2(new_n206), .ZN(new_n208));
  XNOR2_X1  g022(.A(G119), .B(G128), .ZN(new_n209));
  XOR2_X1   g023(.A(KEYINPUT24), .B(G110), .Z(new_n210));
  AOI22_X1  g024(.A1(new_n208), .A2(G110), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n202), .A2(new_n211), .ZN(new_n212));
  OAI22_X1  g026(.A1(new_n208), .A2(G110), .B1(new_n209), .B2(new_n210), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n191), .A2(new_n193), .A3(new_n199), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(new_n201), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT22), .B(G137), .ZN(new_n216));
  INV_X1    g030(.A(G953), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(G221), .A3(G234), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n216), .A2(new_n219), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND4_X1  g036(.A1(new_n212), .A2(KEYINPUT72), .A3(new_n215), .A4(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n212), .A2(new_n215), .A3(new_n222), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT72), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n222), .A2(KEYINPUT71), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT71), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n228), .B1(new_n220), .B2(new_n221), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n230), .B1(new_n212), .B2(new_n215), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n223), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT25), .B1(new_n232), .B2(new_n188), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n189), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n189), .A2(G902), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(G472), .A2(G902), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT32), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT67), .ZN(new_n245));
  INV_X1    g059(.A(G116), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n245), .B1(new_n246), .B2(G119), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n204), .A2(KEYINPUT67), .A3(G116), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(G119), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(new_n248), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT2), .B(G113), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT65), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n253), .B1(new_n199), .B2(G143), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n255), .A2(KEYINPUT65), .A3(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n199), .A2(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT0), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(new_n206), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT64), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n262), .B1(KEYINPUT0), .B2(G128), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n206), .A3(KEYINPUT64), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT66), .B1(new_n255), .B2(G146), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT66), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n199), .A3(G143), .ZN(new_n268));
  AOI22_X1  g082(.A1(new_n266), .A2(new_n268), .B1(new_n255), .B2(G146), .ZN(new_n269));
  AOI22_X1  g083(.A1(new_n259), .A2(new_n265), .B1(new_n269), .B2(new_n261), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT11), .ZN(new_n271));
  INV_X1    g085(.A(G134), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n271), .B1(new_n272), .B2(G137), .ZN(new_n273));
  INV_X1    g087(.A(G137), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(KEYINPUT11), .A3(G134), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n272), .A2(G137), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G131), .ZN(new_n278));
  INV_X1    g092(.A(G131), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n273), .A2(new_n275), .A3(new_n279), .A4(new_n276), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n270), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT30), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n255), .A2(G146), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n267), .B1(G143), .B2(new_n199), .ZN(new_n286));
  NOR3_X1   g100(.A1(new_n255), .A2(KEYINPUT66), .A3(G146), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n284), .B(new_n285), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n258), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n289), .B1(new_n254), .B2(new_n256), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n206), .B1(new_n258), .B2(KEYINPUT1), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n288), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n272), .A2(G137), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n274), .A2(G134), .ZN(new_n294));
  OAI21_X1  g108(.A(G131), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n280), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  AND3_X1   g111(.A1(new_n282), .A2(new_n283), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n283), .B1(new_n282), .B2(new_n297), .ZN(new_n299));
  OAI21_X1  g113(.A(new_n252), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g114(.A1(G237), .A2(G953), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G210), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(KEYINPUT27), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT26), .B(G101), .ZN(new_n304));
  XNOR2_X1  g118(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(new_n252), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n282), .A2(new_n306), .A3(new_n297), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n300), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT31), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(KEYINPUT68), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT68), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n308), .A2(new_n311), .A3(KEYINPUT31), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n307), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n282), .A2(new_n297), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT30), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n282), .A2(new_n297), .A3(new_n283), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n314), .B1(new_n318), .B2(new_n252), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT31), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n319), .A2(KEYINPUT69), .A3(new_n320), .A4(new_n305), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n300), .A2(new_n320), .A3(new_n305), .A4(new_n307), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT69), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n306), .B1(new_n282), .B2(new_n297), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT28), .B1(new_n314), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT28), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n307), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n305), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n321), .A2(new_n324), .A3(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n244), .B1(new_n313), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n300), .A2(new_n307), .ZN(new_n333));
  INV_X1    g147(.A(new_n305), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT29), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n326), .A2(new_n305), .A3(new_n328), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n326), .A2(KEYINPUT29), .A3(new_n305), .A4(new_n328), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n188), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G472), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n332), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n322), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n329), .B1(new_n343), .B2(KEYINPUT69), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n344), .A2(new_n324), .A3(new_n310), .A4(new_n312), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT32), .B1(new_n345), .B2(new_n241), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n240), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT73), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n321), .A2(new_n324), .A3(new_n330), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n308), .A2(new_n311), .A3(KEYINPUT31), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n311), .B1(new_n308), .B2(KEYINPUT31), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n242), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n332), .B(new_n341), .C1(new_n354), .C2(KEYINPUT32), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT73), .A3(new_n240), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n349), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G221), .ZN(new_n358));
  XNOR2_X1  g172(.A(KEYINPUT9), .B(G234), .ZN(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n358), .B1(new_n360), .B2(new_n188), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n190), .A2(G125), .ZN(new_n362));
  OAI21_X1  g176(.A(G146), .B1(new_n195), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(new_n214), .ZN(new_n364));
  NAND2_X1  g178(.A1(KEYINPUT18), .A2(G131), .ZN(new_n365));
  INV_X1    g179(.A(new_n365), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n301), .A2(G143), .A3(G214), .ZN(new_n367));
  AOI21_X1  g181(.A(G143), .B1(new_n301), .B2(G214), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n366), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n301), .A2(G214), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n255), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n301), .A2(G143), .A3(G214), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n365), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n364), .A2(new_n369), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(KEYINPUT84), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT84), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n364), .A2(new_n369), .A3(new_n373), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g192(.A(KEYINPUT17), .B(G131), .C1(new_n367), .C2(new_n368), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n200), .A2(new_n379), .A3(new_n201), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT87), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n200), .A2(new_n379), .A3(KEYINPUT87), .A4(new_n201), .ZN(new_n383));
  OAI21_X1  g197(.A(G131), .B1(new_n367), .B2(new_n368), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n371), .A2(new_n279), .A3(new_n372), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT17), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n383), .A2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n378), .B1(new_n382), .B2(new_n388), .ZN(new_n389));
  XOR2_X1   g203(.A(G113), .B(G122), .Z(new_n390));
  XOR2_X1   g204(.A(KEYINPUT86), .B(G104), .Z(new_n391));
  XNOR2_X1  g205(.A(new_n390), .B(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT19), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(new_n195), .B2(new_n362), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT19), .ZN(new_n395));
  AOI21_X1  g209(.A(G146), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AND3_X1   g210(.A1(new_n194), .A2(G146), .A3(new_n197), .ZN(new_n397));
  OAI21_X1  g211(.A(KEYINPUT85), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n384), .A2(new_n385), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n191), .A2(new_n193), .A3(KEYINPUT19), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT19), .B1(new_n191), .B2(new_n193), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n199), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n201), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n398), .A2(new_n399), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n392), .B1(new_n375), .B2(new_n377), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n389), .A2(new_n392), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(G475), .A2(G902), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n392), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n380), .A2(new_n381), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n387), .A3(new_n383), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n410), .B1(new_n412), .B2(new_n378), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n378), .A2(new_n410), .A3(new_n405), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT88), .ZN(new_n415));
  NOR3_X1   g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n409), .B1(new_n416), .B2(KEYINPUT20), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT20), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n407), .A2(new_n415), .A3(new_n418), .A4(new_n408), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(G478), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n421), .A2(KEYINPUT15), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NOR3_X1   g237(.A1(new_n359), .A2(new_n187), .A3(G953), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n255), .A2(G128), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n206), .A2(G143), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(new_n272), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n427), .A3(G134), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(KEYINPUT90), .A2(G122), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(KEYINPUT90), .A2(G122), .ZN(new_n434));
  OAI21_X1  g248(.A(G116), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n246), .A2(G122), .ZN(new_n436));
  OR2_X1    g250(.A1(new_n436), .A2(KEYINPUT14), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(KEYINPUT92), .A3(KEYINPUT14), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT92), .B1(new_n436), .B2(KEYINPUT14), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n435), .B(new_n437), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n431), .B1(new_n441), .B2(G107), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT90), .ZN(new_n443));
  INV_X1    g257(.A(G122), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n246), .B1(new_n445), .B2(new_n432), .ZN(new_n446));
  INV_X1    g260(.A(new_n436), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT91), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT91), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n435), .A2(new_n449), .A3(new_n436), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G107), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n442), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT13), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n272), .B1(new_n427), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(new_n456), .B(new_n428), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n448), .A2(G107), .A3(new_n450), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n457), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n425), .B1(new_n454), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n457), .ZN(new_n461));
  AND3_X1   g275(.A1(new_n448), .A2(G107), .A3(new_n450), .ZN(new_n462));
  AOI21_X1  g276(.A(G107), .B1(new_n448), .B2(new_n450), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n442), .A2(new_n453), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n465), .A3(new_n424), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n460), .A2(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n423), .B1(new_n467), .B2(new_n188), .ZN(new_n468));
  AOI211_X1 g282(.A(G902), .B(new_n422), .C1(new_n460), .C2(new_n466), .ZN(new_n469));
  NAND2_X1  g283(.A1(G234), .A2(G237), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(G952), .A3(new_n217), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(G898), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n470), .A2(G902), .A3(G953), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n468), .A2(new_n469), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G475), .ZN(new_n478));
  AND2_X1   g292(.A1(new_n383), .A2(new_n387), .ZN(new_n479));
  AOI22_X1  g293(.A1(new_n479), .A2(new_n411), .B1(new_n377), .B2(new_n375), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n392), .A2(KEYINPUT89), .ZN(new_n481));
  AOI21_X1  g295(.A(G902), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n389), .B1(KEYINPUT89), .B2(new_n392), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n478), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n420), .A2(new_n477), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(G104), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT3), .B1(new_n487), .B2(G107), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT3), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n452), .A3(G104), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n487), .A2(G107), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n488), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n492), .A2(new_n493), .A3(G101), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n270), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n490), .A2(new_n491), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT74), .ZN(new_n498));
  INV_X1    g312(.A(G101), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n488), .ZN(new_n500));
  NAND4_X1  g314(.A1(new_n488), .A2(new_n490), .A3(new_n499), .A4(new_n491), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(KEYINPUT74), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n492), .A2(G101), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(KEYINPUT4), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n292), .A2(KEYINPUT10), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n452), .A2(G104), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n491), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n500), .A2(new_n502), .B1(G101), .B2(new_n509), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n496), .A2(new_n505), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT75), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n269), .A2(new_n512), .A3(new_n285), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n284), .B1(new_n286), .B2(new_n287), .ZN(new_n514));
  INV_X1    g328(.A(new_n291), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT75), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n288), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT10), .B1(new_n518), .B2(new_n510), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n281), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n511), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n500), .B2(new_n502), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n509), .A2(G101), .ZN(new_n525));
  AND2_X1   g339(.A1(new_n501), .A2(KEYINPUT74), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n501), .A2(KEYINPUT74), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI22_X1  g342(.A1(new_n524), .A2(new_n495), .B1(new_n528), .B2(new_n506), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n281), .B1(new_n529), .B2(new_n519), .ZN(new_n530));
  XNOR2_X1  g344(.A(G110), .B(G140), .ZN(new_n531));
  AND2_X1   g345(.A1(new_n217), .A2(G227), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n522), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  NOR3_X1   g349(.A1(new_n529), .A2(new_n519), .A3(new_n281), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT12), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n292), .B1(new_n503), .B2(new_n525), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n538), .B1(new_n510), .B2(new_n518), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n537), .B1(new_n539), .B2(new_n521), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n518), .A2(new_n510), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n259), .A2(new_n515), .B1(new_n269), .B2(new_n285), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n528), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n521), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT12), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n536), .B1(new_n540), .B2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n535), .B1(new_n546), .B2(new_n534), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(KEYINPUT76), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT76), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n549), .B(new_n535), .C1(new_n546), .C2(new_n534), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n548), .A2(G469), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G469), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(new_n188), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n540), .A2(new_n545), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n536), .A2(new_n533), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n522), .A2(new_n530), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n533), .ZN(new_n558));
  AOI21_X1  g372(.A(G902), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n553), .B1(new_n559), .B2(new_n552), .ZN(new_n560));
  AOI211_X1 g374(.A(new_n361), .B(new_n486), .C1(new_n551), .C2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT93), .ZN(new_n562));
  OAI21_X1  g376(.A(G210), .B1(G237), .B2(G902), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n563), .B(KEYINPUT82), .Z(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT81), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n288), .B(new_n192), .C1(new_n290), .C2(new_n291), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(new_n270), .B2(new_n192), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n217), .A2(G224), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n568), .A2(KEYINPUT7), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(KEYINPUT7), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n567), .B(new_n571), .C1(new_n270), .C2(new_n192), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n526), .A2(new_n527), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n494), .B(new_n252), .C1(new_n574), .C2(new_n523), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT5), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(new_n204), .A3(G116), .ZN(new_n577));
  OR2_X1    g391(.A1(new_n577), .A2(KEYINPUT77), .ZN(new_n578));
  INV_X1    g392(.A(G113), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n579), .B1(new_n577), .B2(KEYINPUT77), .ZN(new_n580));
  OAI211_X1 g394(.A(new_n578), .B(new_n580), .C1(new_n576), .C2(new_n250), .ZN(new_n581));
  OR2_X1    g395(.A1(new_n250), .A2(new_n251), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n510), .ZN(new_n584));
  XNOR2_X1  g398(.A(G110), .B(G122), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n575), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(KEYINPUT79), .B(KEYINPUT8), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n585), .B(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n581), .A2(new_n582), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n528), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n584), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(new_n573), .B(new_n586), .C1(new_n592), .C2(KEYINPUT80), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n583), .A2(new_n510), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n528), .A2(new_n590), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n588), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT80), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n566), .B(new_n188), .C1(new_n593), .C2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n575), .A2(new_n584), .ZN(new_n600));
  INV_X1    g414(.A(new_n585), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(KEYINPUT6), .A3(new_n586), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n569), .B(KEYINPUT78), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n568), .B(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT6), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n600), .A2(new_n606), .A3(new_n601), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n603), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n599), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n596), .A2(new_n597), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n592), .A2(KEYINPUT80), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n610), .A2(new_n611), .A3(new_n586), .A4(new_n573), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n566), .B1(new_n612), .B2(new_n188), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n565), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(G214), .B1(G237), .B2(G902), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n188), .B1(new_n593), .B2(new_n598), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT81), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n617), .A2(new_n564), .A3(new_n608), .A4(new_n599), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n614), .A2(new_n615), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(KEYINPUT83), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT83), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n614), .A2(new_n618), .A3(new_n621), .A4(new_n615), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n561), .A2(new_n562), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n622), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n361), .B1(new_n551), .B2(new_n560), .ZN(new_n625));
  INV_X1    g439(.A(new_n486), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT93), .B1(new_n624), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n357), .A2(new_n623), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n629), .B(G101), .ZN(G3));
  OAI21_X1  g444(.A(new_n188), .B1(new_n313), .B2(new_n331), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n631), .A2(G472), .B1(new_n345), .B2(new_n241), .ZN(new_n632));
  AND3_X1   g446(.A1(new_n625), .A2(new_n632), .A3(new_n240), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n619), .A2(KEYINPUT94), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT94), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n614), .A2(new_n618), .A3(new_n635), .A4(new_n615), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n476), .B1(new_n634), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n466), .A2(KEYINPUT96), .ZN(new_n638));
  INV_X1    g452(.A(KEYINPUT96), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n464), .A2(new_n465), .A3(new_n639), .A4(new_n424), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n638), .A2(KEYINPUT33), .A3(new_n460), .A4(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT97), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n424), .B1(new_n464), .B2(new_n465), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT33), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT97), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n645), .A2(new_n646), .A3(new_n640), .A4(new_n638), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n642), .A2(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n466), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n644), .B1(new_n649), .B2(new_n643), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT95), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n467), .A2(KEYINPUT95), .A3(new_n644), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n421), .A2(G902), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n648), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n467), .A2(new_n188), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n421), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n419), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n406), .A2(new_n405), .ZN(new_n661));
  OAI211_X1 g475(.A(KEYINPUT88), .B(new_n661), .C1(new_n480), .C2(new_n410), .ZN(new_n662));
  AOI22_X1  g476(.A1(new_n662), .A2(new_n418), .B1(new_n407), .B2(new_n408), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n485), .B1(new_n660), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n659), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n633), .A2(new_n637), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT34), .B(G104), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G6));
  XNOR2_X1  g483(.A(new_n409), .B(KEYINPUT20), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n485), .B1(new_n468), .B2(new_n469), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n633), .A2(new_n637), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT35), .B(G107), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G9));
  INV_X1    g490(.A(new_n235), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(new_n233), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT36), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n230), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n212), .A2(new_n215), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n680), .B(new_n681), .Z(new_n682));
  AOI22_X1  g496(.A1(new_n678), .A2(new_n189), .B1(new_n237), .B2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(KEYINPUT98), .B1(new_n632), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(G472), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n686), .B1(new_n345), .B2(new_n188), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT98), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n687), .A2(new_n354), .A3(new_n688), .A4(new_n683), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n685), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n628), .A3(new_n623), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT37), .B(G110), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G12));
  NAND2_X1  g507(.A1(new_n634), .A2(new_n636), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n345), .A2(new_n244), .B1(G472), .B2(new_n340), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n241), .B1(new_n313), .B2(new_n331), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(new_n243), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n683), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n217), .A2(G900), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n470), .A2(G902), .ZN(new_n701));
  OR3_X1    g515(.A1(new_n700), .A2(KEYINPUT99), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT99), .B1(new_n700), .B2(new_n701), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n471), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n673), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n694), .A2(new_n698), .A3(new_n625), .A4(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G128), .ZN(G30));
  INV_X1    g522(.A(KEYINPUT101), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n704), .B(KEYINPUT39), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n625), .A2(KEYINPUT40), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(KEYINPUT40), .B1(new_n625), .B2(new_n710), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n713), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(KEYINPUT101), .A3(new_n711), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n319), .A2(new_n334), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n314), .A2(new_n325), .A3(new_n305), .ZN(new_n718));
  OR2_X1    g532(.A1(new_n718), .A2(G902), .ZN(new_n719));
  OAI21_X1  g533(.A(G472), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT100), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n697), .A2(new_n722), .A3(new_n332), .ZN(new_n723));
  INV_X1    g537(.A(new_n664), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n468), .A2(new_n469), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n723), .A2(new_n615), .A3(new_n683), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n614), .A2(new_n618), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(KEYINPUT38), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n714), .A2(new_n716), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G143), .ZN(G45));
  INV_X1    g546(.A(new_n704), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n665), .A2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n694), .A2(new_n698), .A3(new_n625), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G146), .ZN(G48));
  NAND2_X1  g550(.A1(new_n559), .A2(new_n552), .ZN(new_n737));
  AOI22_X1  g551(.A1(new_n554), .A2(new_n555), .B1(new_n557), .B2(new_n533), .ZN(new_n738));
  OAI21_X1  g552(.A(G469), .B1(new_n738), .B2(G902), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n737), .A2(new_n739), .A3(KEYINPUT102), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT102), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n741), .B(G469), .C1(new_n738), .C2(G902), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n361), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n347), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n746), .A2(new_n666), .A3(new_n637), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT41), .B(G113), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G15));
  NAND3_X1  g563(.A1(new_n746), .A2(new_n637), .A3(new_n673), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G116), .ZN(G18));
  AOI21_X1  g565(.A(new_n361), .B1(new_n740), .B2(new_n742), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n694), .A2(new_n698), .A3(new_n626), .A4(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G119), .ZN(G21));
  AND2_X1   g568(.A1(new_n752), .A2(new_n475), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n321), .A2(new_n324), .A3(new_n330), .A4(new_n309), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n241), .ZN(new_n757));
  INV_X1    g571(.A(new_n757), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n687), .A2(new_n239), .A3(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n755), .A2(new_n759), .A3(new_n694), .A4(new_n726), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G122), .ZN(G24));
  NOR3_X1   g575(.A1(new_n687), .A2(new_n683), .A3(new_n758), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n694), .A2(new_n762), .A3(new_n734), .A4(new_n752), .ZN(new_n763));
  XOR2_X1   g577(.A(KEYINPUT103), .B(G125), .Z(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G27));
  INV_X1    g579(.A(KEYINPUT42), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n544), .A2(KEYINPUT12), .ZN(new_n767));
  AOI211_X1 g581(.A(new_n537), .B(new_n521), .C1(new_n541), .C2(new_n543), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n522), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n533), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(G469), .A3(new_n535), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n361), .B1(new_n560), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n615), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n614), .B2(new_n618), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n355), .A2(new_n240), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n734), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n766), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n772), .A2(new_n774), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n239), .B1(new_n695), .B2(new_n697), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n778), .A2(KEYINPUT42), .A3(new_n779), .A4(new_n734), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n777), .A2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G131), .ZN(G33));
  INV_X1    g596(.A(KEYINPUT104), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n775), .B2(new_n705), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n778), .A2(KEYINPUT104), .A3(new_n779), .A4(new_n706), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  NAND2_X1  g601(.A1(new_n631), .A2(G472), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n696), .ZN(new_n789));
  AOI21_X1  g603(.A(KEYINPUT109), .B1(new_n789), .B2(new_n684), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT109), .ZN(new_n791));
  NOR3_X1   g605(.A1(new_n632), .A2(new_n791), .A3(new_n683), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT108), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n664), .A2(KEYINPUT106), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT106), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n420), .A2(new_n796), .A3(new_n485), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n659), .A2(new_n795), .A3(KEYINPUT43), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT107), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT43), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n800), .B1(new_n656), .B2(new_n658), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT107), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n801), .A2(new_n802), .A3(new_n795), .A4(new_n797), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n799), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT43), .B1(new_n659), .B2(new_n724), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n794), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  AOI211_X1 g621(.A(KEYINPUT108), .B(new_n805), .C1(new_n799), .C2(new_n803), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n793), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT44), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n793), .B(KEYINPUT44), .C1(new_n807), .C2(new_n808), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT45), .ZN(new_n813));
  INV_X1    g627(.A(new_n550), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n549), .B1(new_n770), .B2(new_n535), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g630(.A(G469), .B1(new_n547), .B2(new_n813), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n553), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n737), .B1(new_n819), .B2(KEYINPUT46), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n548), .A2(new_n550), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n817), .B1(new_n821), .B2(new_n813), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT46), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n822), .A2(new_n823), .A3(new_n553), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n744), .B(new_n710), .C1(new_n820), .C2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT105), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n819), .A2(KEYINPUT46), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n823), .B1(new_n822), .B2(new_n553), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n827), .A2(new_n828), .A3(new_n737), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT105), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n830), .A3(new_n744), .A4(new_n710), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n826), .A2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n811), .A2(new_n774), .A3(new_n812), .A4(new_n832), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(G137), .ZN(G39));
  XNOR2_X1  g648(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n829), .A2(new_n744), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n835), .B1(new_n829), .B2(new_n744), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n355), .A2(new_n240), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n839), .A2(new_n734), .A3(new_n774), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n837), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(new_n190), .ZN(G42));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n725), .A2(KEYINPUT112), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT112), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n845), .B1(new_n468), .B2(new_n469), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n724), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n665), .A2(new_n848), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n624), .A2(new_n849), .A3(new_n476), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n633), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n629), .A2(new_n691), .A3(new_n851), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n747), .A2(new_n750), .A3(new_n760), .A4(new_n753), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n777), .A2(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT113), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n355), .A2(new_n625), .A3(new_n684), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n484), .A2(new_n733), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n670), .A2(new_n844), .A3(new_n846), .A4(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n774), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n855), .B1(new_n856), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n859), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n698), .A3(KEYINPUT113), .A4(new_n625), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n762), .A2(new_n734), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n860), .A2(new_n862), .B1(new_n863), .B2(new_n778), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n852), .A2(new_n853), .A3(new_n854), .A4(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n560), .A2(new_n771), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n682), .A2(new_n237), .ZN(new_n867));
  AND3_X1   g681(.A1(new_n236), .A2(new_n867), .A3(new_n704), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n866), .A2(new_n744), .A3(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n694), .A2(new_n869), .A3(new_n723), .A4(new_n726), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n707), .A2(new_n870), .A3(new_n735), .A4(new_n763), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n871), .B(KEYINPUT52), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n865), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n864), .A2(new_n781), .A3(new_n786), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n629), .A2(new_n691), .A3(new_n851), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n747), .A2(new_n750), .A3(new_n760), .A4(new_n753), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n707), .A2(new_n735), .A3(new_n763), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n879), .A2(KEYINPUT52), .A3(new_n870), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT52), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n871), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT53), .B1(new_n878), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n843), .B1(new_n874), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n873), .B1(new_n865), .B2(new_n872), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n878), .A2(KEYINPUT53), .A3(new_n883), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(KEYINPUT54), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT51), .ZN(new_n890));
  INV_X1    g704(.A(new_n759), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n805), .B1(new_n799), .B2(new_n803), .ZN(new_n892));
  OR3_X1    g706(.A1(new_n892), .A2(KEYINPUT114), .A3(new_n471), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT114), .B1(new_n892), .B2(new_n471), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n774), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n743), .B(KEYINPUT116), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n361), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(new_n837), .B2(new_n838), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n890), .B1(new_n897), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n752), .A2(new_n774), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n902), .B1(new_n893), .B2(new_n894), .ZN(new_n903));
  NOR4_X1   g717(.A1(new_n902), .A2(new_n471), .A3(new_n723), .A4(new_n239), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n659), .A2(new_n664), .ZN(new_n905));
  AOI22_X1  g719(.A1(new_n903), .A2(new_n762), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT118), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n907), .A2(KEYINPUT50), .ZN(new_n908));
  INV_X1    g722(.A(new_n729), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n773), .B1(new_n907), .B2(KEYINPUT50), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n745), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n908), .B1(new_n895), .B2(new_n911), .ZN(new_n912));
  AND3_X1   g726(.A1(new_n895), .A2(new_n908), .A3(new_n911), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n901), .B(new_n906), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n217), .A2(G952), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n915), .B1(new_n904), .B2(new_n666), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT48), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n903), .A2(new_n917), .A3(new_n779), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n917), .B1(new_n903), .B2(new_n779), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n916), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n895), .A2(new_n694), .A3(new_n752), .ZN(new_n921));
  OR2_X1    g735(.A1(new_n921), .A2(KEYINPUT120), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(KEYINPUT120), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n889), .A2(new_n914), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n906), .B1(new_n913), .B2(new_n912), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT115), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n927), .B1(new_n837), .B2(new_n838), .ZN(new_n928));
  INV_X1    g742(.A(new_n838), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(KEYINPUT115), .A3(new_n836), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n899), .B(KEYINPUT117), .Z(new_n932));
  AOI21_X1  g746(.A(new_n896), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n890), .B1(new_n926), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(KEYINPUT119), .ZN(new_n935));
  INV_X1    g749(.A(KEYINPUT119), .ZN(new_n936));
  OAI211_X1 g750(.A(new_n936), .B(new_n890), .C1(new_n926), .C2(new_n933), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  OAI22_X1  g752(.A1(new_n925), .A2(new_n938), .B1(G952), .B2(G953), .ZN(new_n939));
  INV_X1    g753(.A(new_n659), .ZN(new_n940));
  NOR4_X1   g754(.A1(new_n940), .A2(new_n773), .A3(new_n361), .A4(new_n239), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n796), .B1(new_n420), .B2(new_n485), .ZN(new_n942));
  AOI211_X1 g756(.A(KEYINPUT106), .B(new_n484), .C1(new_n417), .C2(new_n419), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT49), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n941), .B(new_n944), .C1(new_n945), .C2(new_n743), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT111), .Z(new_n947));
  AOI21_X1  g761(.A(new_n723), .B1(new_n945), .B2(new_n743), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n947), .A2(new_n729), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n939), .A2(new_n949), .ZN(G75));
  AOI21_X1  g764(.A(new_n188), .B1(new_n886), .B2(new_n887), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(new_n564), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT56), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n603), .A2(new_n607), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(new_n605), .ZN(new_n955));
  XOR2_X1   g769(.A(KEYINPUT121), .B(KEYINPUT55), .Z(new_n956));
  XNOR2_X1  g770(.A(new_n955), .B(new_n956), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n952), .A2(new_n953), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n957), .B1(new_n952), .B2(new_n953), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n217), .A2(G952), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(G51));
  XNOR2_X1  g775(.A(new_n553), .B(KEYINPUT57), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n885), .A2(new_n888), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(KEYINPUT122), .ZN(new_n964));
  INV_X1    g778(.A(new_n738), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT122), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n885), .A2(new_n888), .A3(new_n966), .A4(new_n962), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n964), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n822), .B(KEYINPUT123), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n951), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n960), .B1(new_n968), .B2(new_n970), .ZN(G54));
  AND2_X1   g785(.A1(KEYINPUT58), .A2(G475), .ZN(new_n972));
  OAI211_X1 g786(.A(G902), .B(new_n972), .C1(new_n874), .C2(new_n884), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n973), .B1(new_n413), .B2(new_n414), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n951), .A2(new_n407), .A3(new_n972), .ZN(new_n975));
  INV_X1    g789(.A(new_n960), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT124), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT124), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n974), .A2(new_n975), .A3(new_n979), .A4(new_n976), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(G60));
  NAND2_X1  g795(.A1(G478), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT59), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n885), .A2(new_n888), .A3(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n648), .A2(new_n654), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  AND2_X1   g800(.A1(new_n984), .A2(new_n986), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n984), .A2(new_n986), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n987), .A2(new_n988), .A3(new_n960), .ZN(G63));
  NAND2_X1  g803(.A1(G217), .A2(G902), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT60), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n991), .B1(new_n886), .B2(new_n887), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(new_n682), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT61), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n976), .B1(new_n992), .B2(new_n232), .ZN(new_n997));
  OR3_X1    g811(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n996), .B1(new_n995), .B2(new_n997), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(new_n999), .ZN(G66));
  AOI21_X1  g814(.A(new_n217), .B1(new_n473), .B2(G224), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n852), .A2(new_n853), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1001), .B1(new_n1002), .B2(new_n217), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n954), .B1(G898), .B2(new_n217), .ZN(new_n1004));
  XOR2_X1   g818(.A(new_n1003), .B(new_n1004), .Z(G69));
  AOI21_X1  g819(.A(new_n217), .B1(G227), .B2(G900), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n400), .A2(new_n401), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n318), .B(new_n1007), .ZN(new_n1008));
  INV_X1    g822(.A(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n774), .ZN(new_n1010));
  OR2_X1    g824(.A1(new_n790), .A2(new_n792), .ZN(new_n1011));
  INV_X1    g825(.A(new_n803), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n802), .B1(new_n944), .B2(new_n801), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n806), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1014), .A2(KEYINPUT108), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n892), .A2(new_n794), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1011), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1010), .B1(new_n1017), .B2(KEYINPUT44), .ZN(new_n1018));
  AOI22_X1  g832(.A1(new_n809), .A2(new_n810), .B1(new_n826), .B2(new_n831), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n841), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n694), .A2(new_n779), .A3(new_n726), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1021), .B1(new_n826), .B2(new_n831), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n879), .A2(new_n781), .A3(new_n786), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(G953), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1009), .B1(new_n1025), .B2(new_n699), .ZN(new_n1026));
  INV_X1    g840(.A(KEYINPUT126), .ZN(new_n1027));
  AOI21_X1  g841(.A(new_n1006), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(KEYINPUT125), .ZN(new_n1029));
  INV_X1    g843(.A(new_n841), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n833), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n625), .A2(new_n710), .ZN(new_n1032));
  NOR3_X1   g846(.A1(new_n849), .A2(new_n1032), .A3(new_n1010), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n357), .ZN(new_n1034));
  AND3_X1   g848(.A1(new_n731), .A2(new_n879), .A3(KEYINPUT62), .ZN(new_n1035));
  AOI21_X1  g849(.A(KEYINPUT62), .B1(new_n731), .B2(new_n879), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1034), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n217), .B1(new_n1031), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(new_n1008), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1029), .B1(new_n1026), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g854(.A(new_n1036), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n731), .A2(new_n879), .A3(KEYINPUT62), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1020), .A2(new_n1043), .A3(new_n1034), .ZN(new_n1044));
  AOI21_X1  g858(.A(new_n1009), .B1(new_n1044), .B2(new_n217), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n1045), .A2(KEYINPUT125), .ZN(new_n1046));
  OAI21_X1  g860(.A(new_n1028), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n833), .A2(new_n1024), .A3(new_n1030), .ZN(new_n1048));
  NAND2_X1  g862(.A1(new_n1048), .A2(new_n217), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1008), .B1(new_n1049), .B2(new_n700), .ZN(new_n1050));
  OAI21_X1  g864(.A(KEYINPUT125), .B1(new_n1050), .B2(new_n1045), .ZN(new_n1051));
  INV_X1    g865(.A(new_n1006), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1052), .B1(new_n1050), .B2(KEYINPUT126), .ZN(new_n1053));
  NAND2_X1  g867(.A1(new_n1039), .A2(new_n1029), .ZN(new_n1054));
  NAND3_X1  g868(.A1(new_n1051), .A2(new_n1053), .A3(new_n1054), .ZN(new_n1055));
  AND2_X1   g869(.A1(new_n1047), .A2(new_n1055), .ZN(G72));
  NAND2_X1  g870(.A1(G472), .A2(G902), .ZN(new_n1057));
  XOR2_X1   g871(.A(new_n1057), .B(KEYINPUT63), .Z(new_n1058));
  OAI21_X1  g872(.A(new_n1058), .B1(new_n1044), .B2(new_n1002), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1059), .A2(new_n717), .ZN(new_n1060));
  NAND2_X1  g874(.A1(new_n886), .A2(new_n887), .ZN(new_n1061));
  INV_X1    g875(.A(new_n1058), .ZN(new_n1062));
  AOI21_X1  g876(.A(new_n1062), .B1(new_n335), .B2(new_n308), .ZN(new_n1063));
  AOI21_X1  g877(.A(new_n960), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g878(.A(new_n1058), .B1(new_n1048), .B2(new_n1002), .ZN(new_n1065));
  NAND3_X1  g879(.A1(new_n1065), .A2(new_n334), .A3(new_n319), .ZN(new_n1066));
  NAND3_X1  g880(.A1(new_n1060), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g881(.A(KEYINPUT127), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND4_X1  g883(.A1(new_n1060), .A2(new_n1064), .A3(KEYINPUT127), .A4(new_n1066), .ZN(new_n1070));
  NAND2_X1  g884(.A1(new_n1069), .A2(new_n1070), .ZN(G57));
endmodule


