//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G221), .ZN(new_n188));
  INV_X1    g002(.A(G234), .ZN(new_n189));
  NOR3_X1   g003(.A1(new_n188), .A2(new_n189), .A3(G953), .ZN(new_n190));
  XOR2_X1   g004(.A(new_n187), .B(new_n190), .Z(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G125), .B(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT16), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G125), .ZN(new_n196));
  OR2_X1    g010(.A1(new_n196), .A2(KEYINPUT16), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(G146), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(G146), .B1(new_n194), .B2(new_n197), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G119), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT74), .ZN(new_n203));
  INV_X1    g017(.A(G119), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(G128), .ZN(new_n205));
  NOR3_X1   g019(.A1(new_n201), .A2(KEYINPUT74), .A3(G119), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n202), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  XNOR2_X1  g021(.A(KEYINPUT24), .B(G110), .ZN(new_n208));
  OAI22_X1  g022(.A1(new_n199), .A2(new_n200), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT75), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT23), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(KEYINPUT75), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n211), .A2(new_n213), .A3(G119), .A4(new_n201), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n204), .A2(G128), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n202), .A2(new_n215), .A3(new_n210), .A4(KEYINPUT23), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT76), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT76), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n214), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(G110), .A3(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT77), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G110), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n224), .B1(new_n217), .B2(KEYINPUT76), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT77), .A3(new_n220), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n193), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n198), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n215), .A2(KEYINPUT74), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n203), .A2(new_n204), .A3(G128), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n231), .A2(new_n232), .B1(G119), .B2(new_n201), .ZN(new_n233));
  INV_X1    g047(.A(new_n208), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(G110), .B1(new_n214), .B2(new_n216), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT78), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n236), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT78), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n207), .A2(new_n208), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n230), .B1(new_n237), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n192), .B1(new_n227), .B2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n200), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n244), .A2(new_n198), .B1(new_n233), .B2(new_n234), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n225), .A2(KEYINPUT77), .A3(new_n220), .ZN(new_n246));
  AOI21_X1  g060(.A(KEYINPUT77), .B1(new_n225), .B2(new_n220), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n237), .A2(new_n241), .ZN(new_n249));
  INV_X1    g063(.A(new_n230), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n251), .A3(new_n191), .ZN(new_n252));
  INV_X1    g066(.A(G902), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n243), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT79), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(KEYINPUT25), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(G217), .B1(new_n189), .B2(G902), .ZN(new_n259));
  XOR2_X1   g073(.A(new_n259), .B(KEYINPUT73), .Z(new_n260));
  NAND4_X1  g074(.A1(new_n243), .A2(new_n252), .A3(new_n253), .A4(new_n256), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n243), .A2(new_n252), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n260), .A2(G902), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(KEYINPUT80), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n264), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT9), .B(G234), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n271), .B(KEYINPUT81), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n188), .B1(new_n272), .B2(new_n253), .ZN(new_n273));
  AND2_X1   g087(.A1(KEYINPUT3), .A2(G107), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT3), .A2(G107), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n274), .B1(G104), .B2(new_n275), .ZN(new_n276));
  OR2_X1    g090(.A1(KEYINPUT3), .A2(G107), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT83), .ZN(new_n278));
  INV_X1    g092(.A(G104), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(KEYINPUT83), .A2(G104), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n277), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G101), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n276), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G107), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n280), .A2(new_n285), .A3(new_n281), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n283), .B1(G104), .B2(G107), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n284), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g103(.A(KEYINPUT64), .B(G143), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT1), .B1(new_n290), .B2(G146), .ZN(new_n291));
  INV_X1    g105(.A(G143), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(G146), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(KEYINPUT64), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT64), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G143), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n297), .A3(G146), .ZN(new_n298));
  AOI22_X1  g112(.A1(new_n291), .A2(G128), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT1), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n298), .A2(new_n300), .A3(G128), .A4(new_n294), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n289), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT10), .ZN(new_n304));
  OAI21_X1  g118(.A(G128), .B1(new_n293), .B2(new_n300), .ZN(new_n305));
  AOI21_X1  g119(.A(G146), .B1(new_n295), .B2(new_n297), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n228), .A2(G143), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n304), .B1(new_n308), .B2(new_n301), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n303), .A2(new_n304), .B1(new_n289), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n276), .A2(new_n282), .ZN(new_n311));
  AND2_X1   g125(.A1(KEYINPUT84), .A2(G101), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(KEYINPUT4), .A3(new_n312), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n284), .A2(KEYINPUT4), .ZN(new_n314));
  AND2_X1   g128(.A1(new_n311), .A2(new_n312), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n313), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT68), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT65), .ZN(new_n318));
  AND2_X1   g132(.A1(KEYINPUT0), .A2(G128), .ZN(new_n319));
  NOR2_X1   g133(.A1(KEYINPUT0), .A2(G128), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n318), .B(new_n321), .C1(new_n306), .C2(new_n307), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n298), .A2(new_n319), .A3(new_n294), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n307), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n290), .B2(G146), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n318), .B1(new_n326), .B2(new_n321), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n317), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n295), .A2(new_n297), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n307), .B1(new_n329), .B2(new_n228), .ZN(new_n330));
  INV_X1    g144(.A(new_n321), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT65), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n332), .A2(KEYINPUT68), .A3(new_n323), .A4(new_n322), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n316), .A2(new_n328), .A3(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT11), .ZN(new_n335));
  INV_X1    g149(.A(G134), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n335), .B1(new_n336), .B2(G137), .ZN(new_n337));
  INV_X1    g151(.A(G137), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(KEYINPUT11), .A3(G134), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n336), .A2(G137), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(G131), .ZN(new_n342));
  INV_X1    g156(.A(G131), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n337), .A2(new_n339), .A3(new_n343), .A4(new_n340), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT66), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n344), .A2(new_n345), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n342), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT69), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n339), .A2(new_n340), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n351), .A2(KEYINPUT66), .A3(new_n343), .A4(new_n337), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n344), .A2(new_n345), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(KEYINPUT69), .A3(new_n342), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n310), .A2(new_n334), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(G110), .B(G140), .ZN(new_n358));
  INV_X1    g172(.A(G953), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n359), .A2(G227), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n358), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n356), .B1(new_n310), .B2(new_n334), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AOI221_X4 g179(.A(new_n349), .B1(G131), .B2(new_n341), .C1(new_n352), .C2(new_n353), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT69), .B1(new_n354), .B2(new_n342), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n284), .A2(new_n288), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n369), .A2(new_n308), .A3(new_n301), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n303), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(KEYINPUT12), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n352), .A2(new_n353), .B1(G131), .B2(new_n341), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT12), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n357), .B1(new_n372), .B2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n361), .B(KEYINPUT82), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n365), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(G469), .B1(new_n379), .B2(G902), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n310), .A2(new_n356), .A3(new_n334), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n361), .B1(new_n381), .B2(new_n364), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n357), .B(new_n362), .C1(new_n372), .C2(new_n376), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G469), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(new_n253), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n273), .B1(new_n380), .B2(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(G475), .A2(G902), .ZN(new_n388));
  INV_X1    g202(.A(G237), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n389), .A2(new_n359), .A3(G143), .A4(G214), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n359), .A3(G214), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n390), .B1(new_n392), .B2(new_n329), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G131), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT17), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n290), .A2(new_n391), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n343), .A3(new_n390), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n393), .A2(KEYINPUT17), .A3(G131), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n398), .A2(new_n244), .A3(new_n198), .A4(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n193), .B(G146), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n393), .A2(KEYINPUT91), .ZN(new_n402));
  NAND2_X1  g216(.A1(KEYINPUT18), .A2(G131), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n403), .B1(new_n393), .B2(KEYINPUT90), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT90), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT91), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n396), .A2(new_n406), .A3(new_n407), .A4(new_n390), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G113), .B(G122), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(new_n279), .ZN(new_n412));
  AND3_X1   g226(.A1(new_n400), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n394), .A2(new_n397), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT92), .ZN(new_n415));
  INV_X1    g229(.A(G125), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G140), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n196), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT19), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n193), .A2(KEYINPUT19), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n415), .B1(new_n422), .B2(new_n228), .ZN(new_n423));
  AOI211_X1 g237(.A(KEYINPUT92), .B(G146), .C1(new_n420), .C2(new_n421), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n198), .B(new_n414), .C1(new_n423), .C2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n412), .B1(new_n425), .B2(new_n410), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n388), .B1(new_n413), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT20), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n400), .A2(new_n410), .A3(new_n412), .ZN(new_n429));
  OR2_X1    g243(.A1(new_n423), .A2(new_n424), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n199), .B1(new_n394), .B2(new_n397), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n430), .A2(new_n431), .B1(new_n409), .B2(new_n404), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n429), .B1(new_n432), .B2(new_n412), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(new_n388), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n412), .B1(new_n400), .B2(new_n410), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n253), .B1(new_n413), .B2(new_n436), .ZN(new_n437));
  AOI22_X1  g251(.A1(new_n428), .A2(new_n435), .B1(G475), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n295), .A2(new_n297), .A3(G128), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n201), .A2(G143), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(KEYINPUT13), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT13), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n290), .A2(new_n443), .A3(G128), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n442), .A2(G134), .A3(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT93), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n442), .A2(KEYINPUT93), .A3(G134), .A4(new_n444), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G122), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G116), .ZN(new_n451));
  INV_X1    g265(.A(G116), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G122), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G107), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n453), .A3(new_n285), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n440), .A2(new_n336), .A3(new_n441), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n449), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n450), .A2(G116), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n285), .B1(new_n462), .B2(KEYINPUT14), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT94), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT14), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n451), .A2(new_n453), .A3(new_n465), .ZN(new_n466));
  AND3_X1   g280(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n464), .B1(new_n463), .B2(new_n466), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n440), .A2(new_n336), .A3(new_n441), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n336), .B1(new_n440), .B2(new_n441), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n456), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n272), .A2(G217), .A3(new_n359), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n461), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n459), .B1(new_n447), .B2(new_n448), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n469), .A2(new_n472), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n476), .A2(new_n479), .A3(KEYINPUT95), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT95), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n481), .B(new_n474), .C1(new_n477), .C2(new_n478), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n480), .A2(new_n253), .A3(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(G478), .ZN(new_n484));
  NOR2_X1   g298(.A1(new_n484), .A2(KEYINPUT15), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n485), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n480), .A2(new_n253), .A3(new_n482), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(G952), .ZN(new_n490));
  AOI211_X1 g304(.A(G953), .B(new_n490), .C1(G234), .C2(G237), .ZN(new_n491));
  OAI211_X1 g305(.A(G902), .B(G953), .C1(new_n189), .C2(new_n389), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT96), .ZN(new_n493));
  XNOR2_X1  g307(.A(KEYINPUT21), .B(G898), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n439), .A2(new_n489), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G210), .B1(G237), .B2(G902), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND4_X1  g312(.A1(new_n332), .A2(G125), .A3(new_n323), .A4(new_n322), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n308), .A2(new_n301), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(new_n416), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT86), .B(G224), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(new_n359), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n504), .B(KEYINPUT87), .Z(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n502), .B(new_n506), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT2), .B(G113), .Z(new_n508));
  XNOR2_X1  g322(.A(G116), .B(G119), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n284), .A2(KEYINPUT4), .B1(new_n311), .B2(new_n312), .ZN(new_n511));
  AND3_X1   g325(.A1(new_n311), .A2(KEYINPUT4), .A3(new_n312), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n204), .A2(G116), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n452), .A2(G119), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n514), .A2(new_n515), .A3(KEYINPUT5), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n452), .A2(G119), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n516), .A2(new_n519), .A3(G113), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n508), .A2(new_n509), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n284), .A2(new_n520), .A3(new_n521), .A4(new_n288), .ZN(new_n522));
  XNOR2_X1  g336(.A(G110), .B(G122), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n513), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT6), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n513), .A2(new_n522), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n523), .B(KEYINPUT85), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n526), .A2(KEYINPUT6), .A3(new_n527), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n507), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n523), .B(KEYINPUT8), .Z(new_n532));
  NAND2_X1  g346(.A1(new_n520), .A2(new_n521), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n369), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n532), .B1(new_n534), .B2(new_n522), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT88), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  AOI211_X1 g351(.A(KEYINPUT88), .B(new_n532), .C1(new_n534), .C2(new_n522), .ZN(new_n538));
  INV_X1    g352(.A(new_n502), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n504), .A2(KEYINPUT89), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n504), .A2(KEYINPUT89), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(KEYINPUT7), .A3(new_n541), .ZN(new_n542));
  OAI22_X1  g356(.A1(new_n537), .A2(new_n538), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n504), .A2(KEYINPUT7), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n499), .A2(new_n501), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n524), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n253), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n498), .B1(new_n531), .B2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n502), .B(new_n505), .ZN(new_n549));
  AOI22_X1  g363(.A1(new_n524), .A2(KEYINPUT6), .B1(new_n526), .B2(new_n527), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n526), .A2(KEYINPUT6), .A3(new_n527), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n542), .B1(new_n499), .B2(new_n501), .ZN(new_n553));
  INV_X1    g367(.A(new_n532), .ZN(new_n554));
  INV_X1    g368(.A(new_n522), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n284), .A2(new_n288), .B1(new_n520), .B2(new_n521), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n554), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT88), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n535), .A2(new_n536), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n553), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n524), .A2(new_n545), .ZN(new_n561));
  AOI21_X1  g375(.A(G902), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n552), .A2(new_n562), .A3(new_n497), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n548), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G214), .B1(G237), .B2(G902), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n387), .A2(new_n496), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g382(.A(KEYINPUT26), .B(G101), .ZN(new_n569));
  INV_X1    g383(.A(G210), .ZN(new_n570));
  NOR3_X1   g384(.A1(new_n570), .A2(G237), .A3(G953), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n569), .B(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n573));
  XNOR2_X1  g387(.A(new_n572), .B(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT28), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n350), .A2(new_n328), .A3(new_n333), .A4(new_n355), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n336), .A2(G137), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n338), .A2(G134), .ZN(new_n579));
  OAI21_X1  g393(.A(G131), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT67), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(KEYINPUT67), .B(G131), .C1(new_n578), .C2(new_n579), .ZN(new_n583));
  AOI22_X1  g397(.A1(new_n308), .A2(new_n301), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n510), .B1(new_n584), .B2(new_n354), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n577), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n582), .A2(new_n583), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n354), .A2(new_n500), .A3(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n332), .A2(new_n323), .A3(new_n322), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n588), .B1(new_n589), .B2(new_n373), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n590), .A2(new_n510), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n576), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(KEYINPUT28), .B1(new_n577), .B2(new_n585), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n575), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n575), .B1(new_n577), .B2(new_n585), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n588), .A2(KEYINPUT30), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n328), .A2(new_n333), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n596), .B1(new_n597), .B2(new_n368), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n324), .A2(new_n327), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n599), .A2(new_n348), .B1(new_n354), .B2(new_n584), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n510), .B1(new_n600), .B2(KEYINPUT30), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n595), .B1(new_n598), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT31), .ZN(new_n603));
  INV_X1    g417(.A(new_n596), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n577), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n510), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT30), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n606), .B1(new_n590), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT31), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n610), .A3(new_n595), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n594), .A2(new_n603), .A3(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(G472), .A2(G902), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT71), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT32), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n612), .A2(KEYINPUT71), .A3(new_n613), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT72), .ZN(new_n620));
  INV_X1    g434(.A(new_n613), .ZN(new_n621));
  INV_X1    g435(.A(new_n611), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n610), .B1(new_n609), .B2(new_n595), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n621), .B1(new_n624), .B2(new_n594), .ZN(new_n625));
  INV_X1    g439(.A(new_n586), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n606), .B1(new_n577), .B2(new_n588), .ZN(new_n627));
  OAI21_X1  g441(.A(KEYINPUT28), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n593), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT29), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n575), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n628), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n592), .A2(new_n593), .A3(new_n575), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n605), .A2(new_n608), .B1(new_n577), .B2(new_n585), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n630), .B1(new_n634), .B2(new_n574), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n632), .B(new_n253), .C1(new_n633), .C2(new_n635), .ZN(new_n636));
  AOI22_X1  g450(.A1(new_n625), .A2(KEYINPUT32), .B1(new_n636), .B2(G472), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n619), .A2(new_n620), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n620), .B1(new_n619), .B2(new_n637), .ZN(new_n639));
  OAI211_X1 g453(.A(new_n270), .B(new_n568), .C1(new_n638), .C2(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT97), .B(G101), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G3));
  NAND2_X1  g456(.A1(G469), .A2(G902), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n377), .A2(new_n378), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(new_n364), .B2(new_n363), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n386), .B(new_n643), .C1(new_n385), .C2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n273), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n646), .A2(new_n270), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n616), .A2(new_n618), .ZN(new_n649));
  INV_X1    g463(.A(G472), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n650), .B1(new_n612), .B2(new_n253), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n648), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(new_n495), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT33), .ZN(new_n654));
  OAI211_X1 g468(.A(KEYINPUT99), .B(new_n474), .C1(new_n477), .C2(new_n478), .ZN(new_n655));
  AND2_X1   g469(.A1(new_n476), .A2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT99), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n479), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n654), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g473(.A(KEYINPUT33), .B1(new_n480), .B2(new_n482), .ZN(new_n660));
  OAI211_X1 g474(.A(G478), .B(new_n253), .C1(new_n659), .C2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT100), .B(G478), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n483), .A2(new_n662), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n438), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n552), .A2(new_n562), .A3(KEYINPUT98), .A4(new_n497), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n665), .A2(new_n565), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT98), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n548), .A2(new_n667), .A3(new_n563), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n652), .A2(new_n653), .A3(new_n664), .A4(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT34), .B(G104), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G6));
  INV_X1    g486(.A(new_n489), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n439), .A2(new_n673), .A3(new_n495), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n652), .A2(new_n669), .A3(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT35), .B(G107), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G9));
  NOR2_X1   g491(.A1(new_n649), .A2(new_n651), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n248), .A2(new_n251), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n192), .A2(KEYINPUT36), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n267), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n262), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(KEYINPUT101), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT101), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n262), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n568), .A2(new_n678), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT37), .B(G110), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n688), .B(new_n689), .ZN(G12));
  AND3_X1   g504(.A1(new_n612), .A2(KEYINPUT71), .A3(new_n613), .ZN(new_n691));
  AOI21_X1  g505(.A(KEYINPUT71), .B1(new_n612), .B2(new_n613), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n691), .A2(new_n692), .A3(KEYINPUT32), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n636), .A2(G472), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n694), .B1(new_n617), .B2(new_n614), .ZN(new_n695));
  OAI21_X1  g509(.A(KEYINPUT72), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n619), .A2(new_n637), .A3(new_n620), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n428), .A2(new_n435), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n437), .A2(G475), .ZN(new_n700));
  INV_X1    g514(.A(G900), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n491), .B1(new_n493), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n699), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n673), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n646), .A2(new_n647), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n262), .A2(new_n685), .A3(new_n682), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n685), .B1(new_n262), .B2(new_n682), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n698), .A2(new_n669), .A3(new_n705), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G128), .ZN(G30));
  NOR2_X1   g526(.A1(new_n626), .A2(new_n627), .ZN(new_n713));
  AOI21_X1  g527(.A(G902), .B1(new_n713), .B2(new_n575), .ZN(new_n714));
  INV_X1    g528(.A(new_n634), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n574), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  OAI221_X1 g531(.A(new_n619), .B1(new_n617), .B2(new_n614), .C1(new_n650), .C2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(KEYINPUT102), .ZN(new_n719));
  XOR2_X1   g533(.A(new_n702), .B(KEYINPUT39), .Z(new_n720));
  NAND2_X1  g534(.A1(new_n387), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n721), .A2(new_n722), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n564), .B(KEYINPUT38), .Z(new_n725));
  AOI22_X1  g539(.A1(new_n699), .A2(new_n700), .B1(new_n486), .B2(new_n488), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n709), .A2(new_n565), .A3(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n724), .A2(new_n725), .A3(new_n727), .ZN(new_n728));
  OR3_X1    g542(.A1(new_n719), .A2(new_n723), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n329), .ZN(G45));
  AOI211_X1 g544(.A(new_n702), .B(new_n438), .C1(new_n661), .C2(new_n663), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n698), .A2(new_n669), .A3(new_n710), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(KEYINPUT104), .B(G146), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n732), .B(new_n733), .ZN(G48));
  AOI21_X1  g548(.A(new_n385), .B1(new_n384), .B2(new_n253), .ZN(new_n735));
  AOI211_X1 g549(.A(G469), .B(G902), .C1(new_n382), .C2(new_n383), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n737), .A2(KEYINPUT105), .A3(new_n647), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n291), .A2(G128), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n298), .A2(new_n294), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n369), .B1(new_n741), .B2(new_n301), .ZN(new_n742));
  INV_X1    g556(.A(new_n370), .ZN(new_n743));
  OAI211_X1 g557(.A(new_n350), .B(new_n355), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  AOI22_X1  g558(.A1(new_n744), .A2(new_n374), .B1(new_n371), .B2(new_n375), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n363), .A2(new_n745), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n316), .A2(new_n328), .A3(new_n333), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n309), .A2(new_n289), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n748), .B1(new_n742), .B2(KEYINPUT10), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n368), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n362), .B1(new_n750), .B2(new_n357), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n253), .B1(new_n746), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(G469), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n753), .A2(new_n647), .A3(new_n386), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT105), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n738), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n669), .A2(new_n653), .A3(new_n664), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n759), .B(new_n270), .C1(new_n638), .C2(new_n639), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT41), .B(G113), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G15));
  AND4_X1   g576(.A1(new_n669), .A2(new_n738), .A3(new_n756), .A4(new_n674), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n763), .B(new_n270), .C1(new_n638), .C2(new_n639), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G116), .ZN(G18));
  INV_X1    g579(.A(new_n754), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n669), .ZN(new_n767));
  INV_X1    g581(.A(new_n496), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n767), .A2(new_n768), .A3(new_n709), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n769), .B1(new_n638), .B2(new_n639), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G119), .ZN(G21));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT105), .B1(new_n737), .B2(new_n647), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n735), .A2(new_n736), .A3(new_n755), .A4(new_n273), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n628), .A2(new_n629), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n575), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n621), .B1(new_n777), .B2(new_n624), .ZN(new_n778));
  NOR4_X1   g592(.A1(new_n778), .A2(new_n651), .A3(new_n269), .A4(new_n495), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n666), .A2(new_n668), .A3(new_n726), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(KEYINPUT106), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT106), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n666), .A2(new_n668), .A3(new_n726), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n772), .B1(new_n780), .B2(new_n786), .ZN(new_n787));
  INV_X1    g601(.A(new_n651), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n603), .A2(new_n611), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n574), .B1(new_n628), .B2(new_n629), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n613), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n788), .A2(new_n270), .A3(new_n653), .A4(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n757), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(KEYINPUT107), .A3(new_n785), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n787), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G122), .ZN(G24));
  INV_X1    g610(.A(KEYINPUT108), .ZN(new_n797));
  AOI21_X1  g611(.A(G902), .B1(new_n624), .B2(new_n594), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n791), .B1(new_n798), .B2(new_n650), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n797), .B1(new_n799), .B2(new_n709), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n687), .A2(KEYINPUT108), .A3(new_n788), .A4(new_n791), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n767), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n731), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G125), .ZN(G27));
  INV_X1    g619(.A(KEYINPUT42), .ZN(new_n806));
  AND3_X1   g620(.A1(new_n548), .A2(new_n565), .A3(new_n563), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n706), .A2(new_n808), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n270), .B(new_n809), .C1(new_n638), .C2(new_n639), .ZN(new_n810));
  INV_X1    g624(.A(new_n731), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n806), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n387), .A2(new_n731), .A3(new_n807), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n806), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n625), .A2(KEYINPUT32), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n270), .B1(new_n695), .B2(new_n815), .ZN(new_n816));
  AND2_X1   g630(.A1(new_n816), .A2(KEYINPUT109), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(KEYINPUT109), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n814), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n812), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G131), .ZN(G33));
  XNOR2_X1  g635(.A(new_n705), .B(KEYINPUT110), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n698), .A2(new_n270), .A3(new_n809), .A4(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G134), .ZN(G36));
  NAND2_X1  g638(.A1(new_n661), .A2(new_n663), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(new_n438), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT43), .ZN(new_n827));
  OR3_X1    g641(.A1(new_n827), .A2(new_n678), .A3(new_n709), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT44), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n808), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT45), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n385), .B1(new_n645), .B2(new_n831), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n831), .B2(new_n645), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n643), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT46), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n833), .A2(KEYINPUT46), .A3(new_n643), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n836), .A2(new_n386), .A3(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n647), .A3(new_n720), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n830), .B(new_n840), .C1(new_n829), .C2(new_n828), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G137), .ZN(G39));
  NAND2_X1  g656(.A1(new_n838), .A2(new_n647), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT47), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NOR4_X1   g659(.A1(new_n698), .A2(new_n270), .A3(new_n811), .A4(new_n808), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(G140), .ZN(G42));
  NAND2_X1  g662(.A1(new_n766), .A2(new_n807), .ZN(new_n849));
  OR2_X1    g663(.A1(new_n849), .A2(KEYINPUT118), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(KEYINPUT118), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n850), .A2(new_n491), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n719), .A2(new_n270), .A3(new_n852), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n853), .B(KEYINPUT120), .Z(new_n854));
  NAND4_X1  g668(.A1(new_n854), .A2(new_n438), .A3(new_n663), .A4(new_n661), .ZN(new_n855));
  INV_X1    g669(.A(new_n491), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n827), .A2(new_n269), .A3(new_n856), .A4(new_n799), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n753), .A2(new_n386), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n858), .A2(new_n647), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n807), .B(new_n857), .C1(new_n845), .C2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n827), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n852), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g676(.A(new_n862), .B(KEYINPUT119), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n802), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n725), .A2(new_n565), .A3(new_n754), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n857), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT50), .Z(new_n867));
  NAND4_X1  g681(.A1(new_n855), .A2(new_n860), .A3(new_n864), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT51), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n817), .A2(new_n818), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n863), .A2(new_n873), .ZN(new_n874));
  OR3_X1    g688(.A1(new_n874), .A2(KEYINPUT121), .A3(KEYINPUT48), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n874), .A2(KEYINPUT48), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT122), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n874), .A2(KEYINPUT122), .A3(KEYINPUT48), .ZN(new_n879));
  OAI21_X1  g693(.A(KEYINPUT121), .B1(new_n874), .B2(KEYINPUT48), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n875), .A2(new_n878), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n857), .A2(new_n803), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n882), .A2(G952), .A3(new_n359), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n854), .B2(new_n664), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n870), .A2(new_n871), .A3(new_n881), .A4(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(new_n648), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n678), .A2(new_n886), .A3(new_n653), .A4(new_n567), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n489), .B(KEYINPUT114), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n438), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n688), .B1(new_n887), .B2(new_n889), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n652), .A2(new_n653), .A3(new_n567), .A4(new_n664), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n640), .A2(new_n891), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n890), .B1(new_n892), .B2(KEYINPUT113), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n813), .B1(new_n800), .B2(new_n801), .ZN(new_n894));
  INV_X1    g708(.A(new_n704), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n807), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT115), .B1(new_n896), .B2(new_n888), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT114), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n489), .B(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT115), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n899), .A2(new_n807), .A3(new_n900), .A4(new_n895), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n710), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n894), .B1(new_n902), .B2(new_n698), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n903), .A2(new_n823), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT113), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n640), .A2(new_n905), .A3(new_n891), .ZN(new_n906));
  AND4_X1   g720(.A1(new_n820), .A2(new_n893), .A3(new_n904), .A4(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT107), .B1(new_n793), .B2(new_n785), .ZN(new_n908));
  AND4_X1   g722(.A1(KEYINPUT107), .A2(new_n775), .A3(new_n785), .A4(new_n779), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n764), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n760), .A2(new_n770), .ZN(new_n911));
  OAI21_X1  g725(.A(KEYINPUT112), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n269), .B1(new_n696), .B2(new_n697), .ZN(new_n913));
  AOI22_X1  g727(.A1(new_n913), .A2(new_n759), .B1(new_n698), .B2(new_n769), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT112), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n914), .A2(new_n795), .A3(new_n915), .A4(new_n764), .ZN(new_n916));
  AND2_X1   g730(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n907), .A2(new_n917), .A3(KEYINPUT116), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT116), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n820), .A2(new_n893), .A3(new_n904), .A4(new_n906), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n912), .A2(new_n916), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n919), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n706), .A2(new_n683), .A3(new_n702), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n718), .A2(new_n785), .A3(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n732), .A2(new_n711), .A3(new_n804), .A4(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT52), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n925), .A2(new_n926), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n918), .A2(new_n922), .A3(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT53), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT117), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n929), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n927), .A2(KEYINPUT117), .A3(new_n928), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR4_X1   g749(.A1(new_n920), .A2(new_n931), .A3(new_n911), .A4(new_n910), .ZN(new_n936));
  AOI22_X1  g750(.A1(new_n930), .A2(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT54), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n930), .A2(KEYINPUT53), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT53), .B1(new_n933), .B2(new_n934), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n918), .A2(new_n922), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n940), .B(KEYINPUT54), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n939), .A2(new_n944), .ZN(new_n945));
  OAI22_X1  g759(.A1(new_n885), .A2(new_n945), .B1(G952), .B2(G953), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n270), .A2(new_n647), .A3(new_n565), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT111), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n858), .B(KEYINPUT49), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n725), .A2(new_n949), .A3(new_n826), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n719), .A2(new_n948), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n946), .A2(new_n951), .ZN(G75));
  NOR2_X1   g766(.A1(new_n359), .A2(G952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT56), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n930), .A2(new_n931), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n935), .A2(new_n936), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(G902), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n954), .B1(new_n958), .B2(new_n570), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n550), .A2(new_n551), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(new_n549), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT55), .Z(new_n962));
  AOI21_X1  g776(.A(new_n953), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n962), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n954), .B(new_n964), .C1(new_n958), .C2(new_n570), .ZN(new_n965));
  AND2_X1   g779(.A1(new_n963), .A2(new_n965), .ZN(G51));
  NAND2_X1  g780(.A1(new_n957), .A2(KEYINPUT54), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n939), .ZN(new_n968));
  INV_X1    g782(.A(new_n968), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n643), .B(KEYINPUT57), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n384), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n958), .A2(new_n833), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n953), .B1(new_n971), .B2(new_n972), .ZN(G54));
  INV_X1    g787(.A(new_n958), .ZN(new_n974));
  AND2_X1   g788(.A1(KEYINPUT58), .A2(G475), .ZN(new_n975));
  AND3_X1   g789(.A1(new_n974), .A2(new_n433), .A3(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n433), .B1(new_n974), .B2(new_n975), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n976), .A2(new_n977), .A3(new_n953), .ZN(G60));
  INV_X1    g792(.A(new_n953), .ZN(new_n979));
  NAND2_X1  g793(.A1(G478), .A2(G902), .ZN(new_n980));
  XOR2_X1   g794(.A(new_n980), .B(KEYINPUT59), .Z(new_n981));
  AOI21_X1  g795(.A(new_n981), .B1(new_n939), .B2(new_n944), .ZN(new_n982));
  INV_X1    g796(.A(new_n659), .ZN(new_n983));
  INV_X1    g797(.A(new_n660), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n979), .B1(new_n982), .B2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n968), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(KEYINPUT123), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT123), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n968), .A2(new_n990), .A3(new_n987), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n986), .B1(new_n989), .B2(new_n991), .ZN(G63));
  NAND2_X1  g806(.A1(G217), .A2(G902), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT60), .ZN(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n957), .A2(new_n681), .A3(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT124), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT61), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(KEYINPUT125), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n994), .B1(new_n955), .B2(new_n956), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n979), .B(new_n1000), .C1(new_n1001), .C2(new_n264), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n1001), .A2(KEYINPUT124), .A3(new_n681), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n998), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n263), .B1(new_n937), .B2(new_n994), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1005), .A2(new_n979), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1006), .A2(KEYINPUT125), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1005), .A2(new_n996), .A3(new_n979), .A4(new_n1000), .ZN(new_n1008));
  AOI22_X1  g822(.A1(new_n1004), .A2(new_n1007), .B1(KEYINPUT61), .B2(new_n1008), .ZN(G66));
  INV_X1    g823(.A(new_n503), .ZN(new_n1010));
  OAI21_X1  g824(.A(G953), .B1(new_n1010), .B2(new_n494), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n893), .A2(new_n906), .ZN(new_n1012));
  OR2_X1    g826(.A1(new_n921), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1011), .B1(new_n1014), .B2(G953), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n960), .B1(G898), .B2(new_n359), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(G69));
  AND2_X1   g831(.A1(new_n711), .A2(new_n804), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n873), .A2(new_n785), .A3(new_n840), .ZN(new_n1019));
  AND4_X1   g833(.A1(new_n732), .A2(new_n847), .A3(new_n1018), .A4(new_n1019), .ZN(new_n1020));
  AND2_X1   g834(.A1(new_n841), .A2(new_n823), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1020), .A2(new_n820), .A3(new_n1021), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1022), .A2(KEYINPUT127), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT127), .ZN(new_n1024));
  NAND4_X1  g838(.A1(new_n1020), .A2(new_n1024), .A3(new_n820), .A4(new_n1021), .ZN(new_n1025));
  NAND3_X1  g839(.A1(new_n1023), .A2(new_n359), .A3(new_n1025), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n605), .B1(KEYINPUT30), .B2(new_n600), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(new_n422), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1028), .B1(G900), .B2(G953), .ZN(new_n1029));
  AOI21_X1  g843(.A(KEYINPUT126), .B1(new_n1026), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n359), .B1(G227), .B2(G900), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n729), .A2(new_n732), .A3(new_n1018), .ZN(new_n1033));
  OR2_X1    g847(.A1(new_n1033), .A2(KEYINPUT62), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1033), .A2(KEYINPUT62), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n721), .A2(new_n808), .ZN(new_n1036));
  NOR2_X1   g850(.A1(new_n899), .A2(new_n439), .ZN(new_n1037));
  OAI211_X1 g851(.A(new_n913), .B(new_n1036), .C1(new_n664), .C2(new_n1037), .ZN(new_n1038));
  AND2_X1   g852(.A1(new_n841), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n1034), .A2(new_n847), .A3(new_n1035), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(new_n359), .ZN(new_n1041));
  AOI22_X1  g855(.A1(new_n1026), .A2(new_n1029), .B1(new_n1041), .B2(new_n1028), .ZN(new_n1042));
  XNOR2_X1  g856(.A(new_n1032), .B(new_n1042), .ZN(G72));
  NOR2_X1   g857(.A1(new_n715), .A2(new_n574), .ZN(new_n1044));
  AND3_X1   g858(.A1(new_n1023), .A2(new_n1014), .A3(new_n1025), .ZN(new_n1045));
  NAND2_X1  g859(.A1(G472), .A2(G902), .ZN(new_n1046));
  XOR2_X1   g860(.A(new_n1046), .B(KEYINPUT63), .Z(new_n1047));
  INV_X1    g861(.A(new_n1047), .ZN(new_n1048));
  OAI21_X1  g862(.A(new_n1044), .B1(new_n1045), .B2(new_n1048), .ZN(new_n1049));
  INV_X1    g863(.A(new_n716), .ZN(new_n1050));
  NOR3_X1   g864(.A1(new_n1050), .A2(new_n1044), .A3(new_n1048), .ZN(new_n1051));
  OAI211_X1 g865(.A(new_n940), .B(new_n1051), .C1(new_n942), .C2(new_n943), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1047), .B1(new_n1040), .B2(new_n1013), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n953), .B1(new_n1053), .B2(new_n1050), .ZN(new_n1054));
  AND3_X1   g868(.A1(new_n1049), .A2(new_n1052), .A3(new_n1054), .ZN(G57));
endmodule


