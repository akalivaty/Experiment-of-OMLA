//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 0 1 0 0 1 0 1 1 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n450, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n528, new_n529, new_n530, new_n531, new_n532, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n542, new_n544,
    new_n545, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n573, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n608, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XOR2_X1   g016(.A(KEYINPUT64), .B(G108), .Z(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT65), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G2104), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n464), .A2(new_n466), .A3(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n462), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT68), .ZN(new_n470));
  NAND2_X1  g045(.A1(G101), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n472), .B1(new_n473), .B2(G137), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n470), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n464), .A2(new_n466), .A3(G137), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n471), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n477), .A2(KEYINPUT68), .A3(new_n462), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n469), .B1(new_n475), .B2(new_n478), .ZN(G160));
  NAND2_X1  g054(.A1(new_n464), .A2(new_n466), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n480), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(new_n462), .B2(G112), .ZN(new_n485));
  NOR2_X1   g060(.A1(G100), .A2(G2105), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n487), .A2(KEYINPUT69), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n487), .A2(KEYINPUT69), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n482), .B(new_n484), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  NAND4_X1  g066(.A1(new_n464), .A2(new_n466), .A3(G138), .A4(new_n462), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n473), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n464), .A2(new_n466), .A3(G126), .A4(G2105), .ZN(new_n496));
  INV_X1    g071(.A(G114), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2105), .ZN(new_n498));
  OAI211_X1 g073(.A(new_n498), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n494), .A2(new_n495), .A3(new_n496), .A4(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(G164));
  XNOR2_X1  g076(.A(KEYINPUT5), .B(G543), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(KEYINPUT5), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(G543), .ZN(new_n512));
  AND2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  OAI211_X1 g089(.A(new_n510), .B(new_n512), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G88), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n507), .A2(new_n508), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n505), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(new_n515), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G89), .ZN(new_n520));
  AND3_X1   g095(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT70), .B(G51), .ZN(new_n522));
  OAI221_X1 g097(.A(new_n520), .B1(KEYINPUT7), .B2(new_n521), .C1(new_n507), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n502), .A2(G63), .ZN(new_n524));
  NAND3_X1  g099(.A1(KEYINPUT7), .A2(G76), .A3(G543), .ZN(new_n525));
  AOI21_X1  g100(.A(new_n504), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n523), .A2(new_n526), .ZN(G168));
  AOI22_X1  g102(.A1(new_n502), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n504), .ZN(new_n529));
  INV_X1    g104(.A(G52), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n507), .A2(new_n530), .B1(new_n515), .B2(new_n531), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n529), .A2(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  AOI22_X1  g109(.A1(new_n502), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n504), .ZN(new_n536));
  INV_X1    g111(.A(G43), .ZN(new_n537));
  INV_X1    g112(.A(G81), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n507), .A2(new_n537), .B1(new_n515), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G860), .ZN(G153));
  AND3_X1   g116(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G36), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n542), .A2(new_n545), .ZN(G188));
  OR2_X1    g121(.A1(KEYINPUT72), .A2(G65), .ZN(new_n547));
  NAND2_X1  g122(.A1(KEYINPUT72), .A2(G65), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n547), .A2(new_n510), .A3(new_n512), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(KEYINPUT73), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT73), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n549), .A2(new_n553), .A3(new_n550), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n552), .A2(G651), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n515), .A2(KEYINPUT71), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT71), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n502), .A2(new_n506), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G91), .ZN(new_n560));
  INV_X1    g135(.A(G53), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT9), .B1(new_n507), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT9), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n506), .A2(new_n563), .A3(G53), .A4(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n555), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT74), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n555), .A2(new_n568), .A3(new_n560), .A4(new_n565), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(G168), .ZN(G286));
  INV_X1    g146(.A(G166), .ZN(G303));
  NAND2_X1  g147(.A1(new_n559), .A2(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(G651), .B1(new_n502), .B2(G74), .ZN(new_n574));
  INV_X1    g149(.A(new_n507), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G49), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n573), .A2(new_n574), .A3(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(new_n559), .A2(G86), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n510), .A2(new_n512), .ZN(new_n580));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(G651), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n575), .A2(G48), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n582), .A2(KEYINPUT75), .A3(G651), .ZN(new_n587));
  NAND4_X1  g162(.A1(new_n578), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(G305));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  XNOR2_X1  g164(.A(KEYINPUT76), .B(G85), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n507), .A2(new_n589), .B1(new_n515), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT77), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n591), .B(new_n592), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n502), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OR2_X1    g169(.A1(new_n594), .A2(new_n504), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n593), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  AOI21_X1  g173(.A(new_n598), .B1(new_n559), .B2(G92), .ZN(new_n599));
  INV_X1    g174(.A(G92), .ZN(new_n600));
  AOI211_X1 g175(.A(KEYINPUT10), .B(new_n600), .C1(new_n556), .C2(new_n558), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n502), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G54), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n602), .A2(new_n504), .B1(new_n603), .B2(new_n507), .ZN(new_n604));
  NOR3_X1   g179(.A1(new_n599), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n597), .B1(new_n605), .B2(G868), .ZN(G284));
  OAI21_X1  g181(.A(new_n597), .B1(new_n605), .B2(G868), .ZN(G321));
  NAND2_X1  g182(.A1(G286), .A2(G868), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT78), .Z(new_n609));
  XNOR2_X1  g184(.A(G299), .B(KEYINPUT79), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G297));
  OAI21_X1  g186(.A(new_n609), .B1(new_n610), .B2(G868), .ZN(G280));
  INV_X1    g187(.A(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n605), .B1(new_n613), .B2(G860), .ZN(G148));
  NAND2_X1  g189(.A1(new_n605), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n616), .B1(G868), .B2(new_n540), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n483), .A2(G2104), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n481), .A2(G123), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT81), .Z(new_n624));
  NAND2_X1  g199(.A1(new_n483), .A2(G135), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT80), .Z(new_n626));
  OR2_X1    g201(.A1(G99), .A2(G2105), .ZN(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n628));
  AND3_X1   g203(.A1(new_n624), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n622), .A2(new_n630), .ZN(G156));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2435), .ZN(new_n633));
  XOR2_X1   g208(.A(G2427), .B(G2438), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n635), .A2(KEYINPUT14), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  AND2_X1   g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n638), .A2(new_n640), .ZN(new_n642));
  XOR2_X1   g217(.A(G2451), .B(G2454), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT82), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  OR3_X1    g221(.A1(new_n641), .A2(new_n642), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n646), .B1(new_n641), .B2(new_n642), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n647), .A2(G14), .A3(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(G401));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  XOR2_X1   g226(.A(G2067), .B(G2678), .Z(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n651), .B1(new_n655), .B2(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(G2096), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2100), .ZN(new_n658));
  AND2_X1   g233(.A1(new_n655), .A2(KEYINPUT17), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n653), .A2(new_n654), .ZN(new_n660));
  AOI21_X1  g235(.A(KEYINPUT18), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n658), .B(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(G227));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  NOR2_X1   g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n665), .ZN(new_n671));
  OR2_X1    g246(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT20), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n667), .A2(new_n669), .A3(new_n671), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n674), .B(new_n675), .C1(new_n673), .C2(new_n672), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT21), .B(G1986), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1991), .B(G1996), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT22), .B(G1981), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n680), .B(new_n681), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(G229));
  XNOR2_X1  g258(.A(KEYINPUT83), .B(G29), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G35), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G162), .B2(new_n685), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n688));
  INV_X1    g263(.A(G2090), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n687), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(G160), .ZN(new_n692));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT24), .B(G34), .Z(new_n694));
  OAI22_X1  g269(.A1(new_n692), .A2(new_n693), .B1(new_n684), .B2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(G2084), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(G5), .A2(G16), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(G171), .B2(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n481), .A2(G129), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n483), .A2(G141), .ZN(new_n701));
  NAND3_X1  g276(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n702));
  XOR2_X1   g277(.A(new_n702), .B(KEYINPUT26), .Z(new_n703));
  NAND3_X1  g278(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n704), .B(KEYINPUT91), .ZN(new_n705));
  NAND4_X1  g280(.A1(new_n700), .A2(new_n701), .A3(new_n703), .A4(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT92), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n706), .A2(new_n707), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G29), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G29), .B2(G32), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT27), .B(G1996), .ZN(new_n714));
  OAI221_X1 g289(.A(new_n697), .B1(G1961), .B2(new_n699), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n715), .B(KEYINPUT94), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n685), .A2(G27), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G164), .B2(new_n685), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(G2078), .Z(new_n719));
  XOR2_X1   g294(.A(KEYINPUT30), .B(G28), .Z(new_n720));
  NOR2_X1   g295(.A1(KEYINPUT31), .A2(G11), .ZN(new_n721));
  AND2_X1   g296(.A1(KEYINPUT31), .A2(G11), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n719), .B1(G29), .B2(new_n720), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  AND2_X1   g298(.A1(new_n699), .A2(G1961), .ZN(new_n724));
  NAND3_X1  g299(.A1(new_n624), .A2(new_n626), .A3(new_n628), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n725), .A2(new_n685), .ZN(new_n726));
  NOR2_X1   g301(.A1(G16), .A2(G21), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G168), .B2(G16), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT93), .B(G1966), .Z(new_n729));
  OAI22_X1  g304(.A1(new_n728), .A2(new_n729), .B1(new_n695), .B2(new_n696), .ZN(new_n730));
  NOR4_X1   g305(.A1(new_n723), .A2(new_n724), .A3(new_n726), .A4(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(G29), .A2(G33), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n473), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  INV_X1    g308(.A(G139), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n473), .A2(new_n462), .ZN(new_n735));
  OAI22_X1  g310(.A1(new_n733), .A2(new_n462), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT25), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n732), .B1(new_n739), .B2(G29), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n728), .A2(new_n729), .B1(G2072), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n713), .A2(new_n714), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n716), .A2(new_n731), .A3(new_n741), .A4(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(G16), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n744), .A2(G4), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n605), .B2(new_n744), .ZN(new_n746));
  INV_X1    g321(.A(G1348), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n685), .A2(G26), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n481), .A2(G128), .ZN(new_n752));
  OR2_X1    g327(.A1(G104), .A2(G2105), .ZN(new_n753));
  OAI211_X1 g328(.A(new_n753), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT88), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n752), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n483), .A2(KEYINPUT87), .A3(G140), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT87), .ZN(new_n760));
  INV_X1    g335(.A(G140), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n735), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n759), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g338(.A1(new_n758), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n751), .B1(new_n764), .B2(new_n693), .ZN(new_n765));
  INV_X1    g340(.A(G2067), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n744), .A2(G19), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(new_n540), .B2(new_n744), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(G1341), .Z(new_n770));
  NAND3_X1  g345(.A1(new_n748), .A2(new_n767), .A3(new_n770), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT90), .Z(new_n772));
  NOR2_X1   g347(.A1(new_n743), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT36), .ZN(new_n774));
  INV_X1    g349(.A(KEYINPUT86), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT85), .ZN(new_n776));
  NOR2_X1   g351(.A1(G288), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(G288), .A2(new_n776), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n744), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NOR2_X1   g355(.A1(G16), .A2(G23), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n775), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  XOR2_X1   g358(.A(KEYINPUT33), .B(G1976), .Z(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NOR3_X1   g360(.A1(new_n780), .A2(new_n775), .A3(new_n781), .ZN(new_n786));
  NOR3_X1   g361(.A1(new_n783), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  OR3_X1    g362(.A1(new_n780), .A2(new_n775), .A3(new_n781), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n784), .B1(new_n788), .B2(new_n782), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n744), .A2(G22), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G166), .B2(new_n744), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(G1971), .Z(new_n793));
  NAND2_X1  g368(.A1(new_n744), .A2(G6), .ZN(new_n794));
  INV_X1    g369(.A(G305), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n794), .B1(new_n795), .B2(new_n744), .ZN(new_n796));
  XOR2_X1   g371(.A(KEYINPUT32), .B(G1981), .Z(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n790), .A2(KEYINPUT34), .A3(new_n793), .A4(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n785), .B1(new_n783), .B2(new_n786), .ZN(new_n800));
  NAND3_X1  g375(.A1(new_n788), .A2(new_n784), .A3(new_n782), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n800), .A2(new_n793), .A3(new_n801), .A4(new_n798), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT34), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n799), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n684), .A2(G25), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n481), .A2(G119), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT84), .Z(new_n808));
  INV_X1    g383(.A(G131), .ZN(new_n809));
  NOR2_X1   g384(.A1(G95), .A2(G2105), .ZN(new_n810));
  OAI21_X1  g385(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n735), .A2(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n808), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n806), .B1(new_n813), .B2(new_n684), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT35), .B(G1991), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n814), .B(new_n815), .Z(new_n816));
  NAND2_X1  g391(.A1(new_n744), .A2(G24), .ZN(new_n817));
  INV_X1    g392(.A(G290), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(new_n744), .ZN(new_n819));
  INV_X1    g394(.A(G1986), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n816), .A2(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n774), .B1(new_n805), .B2(new_n823), .ZN(new_n824));
  AOI211_X1 g399(.A(KEYINPUT36), .B(new_n822), .C1(new_n799), .C2(new_n804), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n691), .B(new_n773), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(G299), .A2(G16), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n744), .A2(KEYINPUT23), .A3(G20), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT23), .ZN(new_n829));
  INV_X1    g404(.A(G20), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(G16), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n827), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT96), .B(G1956), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n832), .B(new_n833), .Z(new_n834));
  NOR2_X1   g409(.A1(new_n740), .A2(G2072), .ZN(new_n835));
  NOR3_X1   g410(.A1(new_n826), .A2(new_n834), .A3(new_n835), .ZN(G311));
  INV_X1    g411(.A(new_n773), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n805), .A2(new_n823), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT36), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n805), .A2(new_n774), .A3(new_n823), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n837), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n834), .ZN(new_n842));
  INV_X1    g417(.A(new_n835), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .A4(new_n691), .ZN(G150));
  NAND2_X1  g419(.A1(new_n605), .A2(G559), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT38), .Z(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT39), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n502), .A2(G67), .ZN(new_n848));
  NAND2_X1  g423(.A1(G80), .A2(G543), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n504), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT97), .ZN(new_n852));
  OAI211_X1 g427(.A(G55), .B(G543), .C1(new_n513), .C2(new_n514), .ZN(new_n853));
  INV_X1    g428(.A(G93), .ZN(new_n854));
  OAI211_X1 g429(.A(new_n852), .B(new_n853), .C1(new_n515), .C2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n502), .A2(new_n506), .A3(G93), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n852), .B1(new_n857), .B2(new_n853), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n851), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT98), .ZN(new_n860));
  INV_X1    g435(.A(new_n540), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT98), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n851), .B(new_n862), .C1(new_n856), .C2(new_n858), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n860), .A2(new_n861), .A3(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n859), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n865), .A2(new_n862), .A3(new_n540), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  XOR2_X1   g442(.A(new_n847), .B(new_n867), .Z(new_n868));
  INV_X1    g443(.A(G860), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(KEYINPUT99), .Z(new_n871));
  NAND2_X1  g446(.A1(new_n859), .A2(G860), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n872), .B(KEYINPUT100), .Z(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(KEYINPUT37), .Z(new_n874));
  NAND2_X1  g449(.A1(new_n871), .A2(new_n874), .ZN(G145));
  NAND2_X1  g450(.A1(new_n496), .A2(new_n499), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT101), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n496), .A2(new_n499), .A3(KEYINPUT101), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n494), .A2(new_n495), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT102), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n764), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(KEYINPUT102), .B1(new_n758), .B2(new_n763), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n883), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n710), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n462), .A2(G118), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT103), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n891), .B(G2104), .C1(G106), .C2(G2105), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n483), .A2(G142), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n481), .A2(G130), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n889), .A2(new_n708), .A3(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n895), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n709), .B2(new_n710), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n885), .A2(new_n886), .A3(new_n883), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n888), .A2(new_n896), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n896), .ZN(new_n901));
  INV_X1    g476(.A(new_n899), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n901), .B1(new_n902), .B2(new_n887), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n739), .ZN(new_n905));
  NAND2_X1  g480(.A1(G160), .A2(new_n490), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(G160), .A2(new_n490), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n629), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n725), .B1(new_n907), .B2(new_n908), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n905), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n910), .A2(new_n905), .A3(new_n911), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n904), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n910), .A2(new_n905), .A3(new_n911), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n900), .B(new_n903), .C1(new_n916), .C2(new_n912), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n813), .B(new_n620), .Z(new_n918));
  AND3_X1   g493(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n918), .B1(new_n915), .B2(new_n917), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(G37), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n923), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g499(.A1(new_n593), .A2(G303), .A3(new_n595), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AOI21_X1  g501(.A(G303), .B1(new_n593), .B2(new_n595), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n779), .B(new_n778), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(G290), .A2(G166), .ZN(new_n929));
  INV_X1    g504(.A(new_n779), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n929), .B(new_n925), .C1(new_n930), .C2(new_n777), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n795), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n928), .A2(new_n931), .A3(new_n795), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g510(.A1(KEYINPUT104), .A2(KEYINPUT42), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n937), .B1(KEYINPUT104), .B2(KEYINPUT42), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n936), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  XOR2_X1   g515(.A(new_n867), .B(new_n615), .Z(new_n941));
  AND3_X1   g516(.A1(new_n567), .A2(new_n605), .A3(new_n569), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n605), .B1(new_n567), .B2(new_n569), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT41), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n946), .B1(new_n942), .B2(new_n943), .ZN(new_n947));
  INV_X1    g522(.A(new_n605), .ZN(new_n948));
  NAND2_X1  g523(.A1(G299), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n567), .A2(new_n605), .A3(new_n569), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(KEYINPUT41), .A3(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n945), .B1(new_n952), .B2(new_n941), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n940), .B(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(G868), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n955), .B1(G868), .B2(new_n865), .ZN(G295));
  OAI21_X1  g531(.A(new_n955), .B1(G868), .B2(new_n865), .ZN(G331));
  INV_X1    g532(.A(KEYINPUT43), .ZN(new_n958));
  AOI21_X1  g533(.A(G301), .B1(G168), .B2(KEYINPUT105), .ZN(new_n959));
  INV_X1    g534(.A(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT105), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n961), .B1(new_n523), .B2(new_n526), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n864), .A2(new_n866), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n864), .B2(new_n866), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n962), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n867), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n864), .A2(new_n866), .A3(new_n962), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n959), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n965), .A2(new_n969), .A3(new_n944), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT106), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n952), .B1(new_n969), .B2(new_n965), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n965), .A2(new_n969), .A3(new_n944), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n971), .B(new_n935), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n965), .A2(new_n969), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n947), .A2(new_n951), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n934), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(new_n932), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n977), .B(new_n970), .C1(new_n979), .C2(KEYINPUT106), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n974), .A2(new_n922), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT107), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT107), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n974), .A2(new_n980), .A3(new_n983), .A4(new_n922), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n958), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n935), .B1(new_n972), .B2(new_n973), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n977), .A2(new_n979), .A3(new_n970), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n986), .A2(new_n922), .A3(new_n987), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n988), .A2(new_n958), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT44), .B1(new_n985), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(KEYINPUT43), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n974), .A2(new_n980), .A3(new_n958), .A4(new_n922), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n990), .B1(KEYINPUT44), .B2(new_n994), .ZN(G397));
  AOI21_X1  g570(.A(G1384), .B1(new_n880), .B2(new_n882), .ZN(new_n996));
  INV_X1    g571(.A(new_n469), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT109), .B(G40), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(KEYINPUT68), .B1(new_n477), .B2(new_n462), .ZN(new_n1000));
  AOI211_X1 g575(.A(new_n470), .B(G2105), .C1(new_n476), .C2(new_n471), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n997), .B(new_n999), .C1(new_n1000), .C2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n996), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n711), .B(G1996), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n764), .B(G2067), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n813), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n815), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n815), .ZN(new_n1010));
  INV_X1    g585(.A(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1007), .A2(new_n1009), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n820), .B2(new_n818), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G290), .A2(G1986), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1004), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G1384), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n500), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1002), .B1(KEYINPUT50), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT50), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n496), .A2(new_n499), .A3(KEYINPUT101), .ZN(new_n1021));
  AOI21_X1  g596(.A(KEYINPUT101), .B1(new_n496), .B2(new_n499), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1020), .B(new_n1017), .C1(new_n1023), .C2(new_n881), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT111), .B1(new_n1025), .B2(G2090), .ZN(new_n1026));
  OAI211_X1 g601(.A(KEYINPUT45), .B(new_n1017), .C1(new_n1023), .C2(new_n881), .ZN(new_n1027));
  AOI211_X1 g602(.A(new_n469), .B(new_n998), .C1(new_n475), .C2(new_n478), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1003), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1018), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(KEYINPUT110), .B(G1971), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1019), .A2(new_n1034), .A3(new_n689), .A4(new_n1024), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1026), .A2(new_n1033), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G303), .A2(G8), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT112), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT55), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(KEYINPUT55), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1037), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(G303), .A2(G8), .A3(new_n1040), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1036), .A2(G8), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G1976), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1045), .B1(new_n778), .B2(new_n779), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT113), .B(G8), .Z(new_n1047));
  INV_X1    g622(.A(new_n996), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(new_n1002), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT52), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1049), .ZN(new_n1051));
  OAI21_X1  g626(.A(G1976), .B1(new_n930), .B2(new_n777), .ZN(new_n1052));
  AOI21_X1  g627(.A(KEYINPUT52), .B1(G288), .B2(new_n1045), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  OR2_X1    g629(.A1(G305), .A2(G1981), .ZN(new_n1055));
  XOR2_X1   g630(.A(KEYINPUT114), .B(G86), .Z(new_n1056));
  OAI211_X1 g631(.A(new_n586), .B(new_n583), .C1(new_n515), .C2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(G1981), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1055), .A2(KEYINPUT49), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1058), .B1(G305), .B2(G1981), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT49), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1059), .A2(new_n1051), .A3(new_n1062), .ZN(new_n1063));
  AND3_X1   g638(.A1(new_n1050), .A2(new_n1054), .A3(new_n1063), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1044), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1028), .B1(KEYINPUT50), .B2(new_n1018), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n996), .A2(new_n1020), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1067), .A2(new_n1068), .A3(G2090), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1069), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1047), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1066), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1065), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(G1966), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1028), .B1(new_n996), .B2(KEYINPUT45), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n500), .A2(new_n1017), .A3(new_n1003), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT115), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT115), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n500), .A2(new_n1079), .A3(new_n1017), .A4(new_n1003), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1075), .B1(new_n1076), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1018), .A2(KEYINPUT50), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1024), .A2(new_n1028), .A3(new_n696), .A4(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT116), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT116), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1019), .A2(new_n1086), .A3(new_n696), .A4(new_n1024), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1082), .A2(new_n1085), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G8), .ZN(new_n1089));
  NOR2_X1   g664(.A1(G168), .A2(new_n1071), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(KEYINPUT121), .A3(KEYINPUT51), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1090), .B1(new_n1088), .B2(G8), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT51), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1094), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1088), .A2(new_n1047), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1090), .A2(KEYINPUT51), .ZN(new_n1099));
  AOI22_X1  g674(.A1(new_n1093), .A2(new_n1097), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1088), .A2(G286), .A3(new_n1047), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT62), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1104));
  AOI21_X1  g679(.A(KEYINPUT121), .B1(new_n1092), .B2(KEYINPUT51), .ZN(new_n1105));
  NOR3_X1   g680(.A1(new_n1095), .A2(new_n1094), .A3(new_n1096), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1104), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT62), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(new_n1108), .A3(new_n1101), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n1031), .A2(G2078), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT53), .ZN(new_n1111));
  INV_X1    g686(.A(G1961), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1110), .A2(new_n1111), .B1(new_n1112), .B2(new_n1025), .ZN(new_n1113));
  OR4_X1    g688(.A1(new_n1111), .A2(new_n1076), .A3(new_n1081), .A4(G2078), .ZN(new_n1114));
  AOI21_X1  g689(.A(G301), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1103), .A2(new_n1109), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1107), .A2(new_n1101), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1025), .A2(new_n747), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1048), .A2(new_n1002), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n766), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1118), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G1956), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1122), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n566), .B(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g700(.A(KEYINPUT56), .B(G2072), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1027), .A2(new_n1028), .A3(new_n1030), .A4(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1123), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1121), .A2(new_n1128), .A3(new_n605), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n566), .B(KEYINPUT57), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1018), .A2(KEYINPUT50), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1131), .A2(new_n1002), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1023), .A2(new_n881), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT50), .B1(new_n1133), .B2(G1384), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1956), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1127), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1130), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  AND2_X1   g712(.A1(new_n1129), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n605), .A2(KEYINPUT60), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1118), .A2(new_n1120), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1139), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1141));
  OAI22_X1  g716(.A1(new_n1140), .A2(new_n1141), .B1(KEYINPUT60), .B2(new_n605), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT119), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1137), .A2(new_n1128), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT61), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  AOI211_X1 g721(.A(KEYINPUT119), .B(KEYINPUT61), .C1(new_n1137), .C2(new_n1128), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1142), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT120), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1149), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1150));
  XNOR2_X1  g725(.A(KEYINPUT58), .B(G1341), .ZN(new_n1151));
  OAI22_X1  g726(.A1(new_n1119), .A2(new_n1151), .B1(new_n1031), .B2(G1996), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n540), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(KEYINPUT59), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1152), .A2(new_n1155), .A3(new_n540), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1154), .A2(new_n1156), .ZN(new_n1157));
  NAND4_X1  g732(.A1(new_n1137), .A2(new_n1128), .A3(KEYINPUT120), .A4(KEYINPUT61), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1150), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(new_n1138), .B1(new_n1148), .B2(new_n1159), .ZN(new_n1160));
  OAI211_X1 g735(.A(new_n1027), .B(G40), .C1(new_n996), .C2(new_n1003), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT123), .B(G2078), .ZN(new_n1162));
  OR3_X1    g737(.A1(new_n1161), .A2(new_n1111), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1113), .B1(new_n692), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(G171), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1113), .A2(G301), .A3(new_n1114), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1165), .A2(KEYINPUT54), .A3(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1168));
  NOR2_X1   g743(.A1(new_n1164), .A2(G171), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1168), .B1(new_n1169), .B2(new_n1115), .ZN(new_n1170));
  NAND4_X1  g745(.A1(new_n1117), .A2(new_n1160), .A3(new_n1167), .A4(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1074), .B1(new_n1116), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(G288), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1063), .A2(new_n1045), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g749(.A(new_n1049), .B1(new_n1174), .B2(new_n1055), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1044), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1175), .B1(new_n1176), .B2(new_n1064), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1088), .A2(G168), .A3(new_n1047), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT117), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n1178), .B(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT63), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1036), .A2(G8), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1181), .B1(new_n1182), .B2(new_n1066), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1065), .A2(new_n1180), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1184), .A2(KEYINPUT118), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT118), .ZN(new_n1186));
  NAND4_X1  g761(.A1(new_n1065), .A2(new_n1180), .A3(new_n1186), .A4(new_n1183), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1185), .A2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g763(.A(KEYINPUT63), .B1(new_n1073), .B2(new_n1180), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1177), .B1(new_n1188), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1016), .B1(new_n1172), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1015), .A2(new_n1004), .ZN(new_n1192));
  XOR2_X1   g767(.A(new_n1192), .B(KEYINPUT48), .Z(new_n1193));
  AOI21_X1  g768(.A(new_n1193), .B1(new_n1012), .B2(new_n1004), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1004), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n764), .A2(new_n766), .ZN(new_n1197));
  AOI21_X1  g772(.A(new_n1195), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  XOR2_X1   g773(.A(new_n1198), .B(KEYINPUT124), .Z(new_n1199));
  INV_X1    g774(.A(KEYINPUT46), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1200), .B1(new_n1195), .B2(G1996), .ZN(new_n1201));
  XNOR2_X1  g776(.A(new_n1201), .B(KEYINPUT125), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1195), .B1(new_n711), .B2(new_n1006), .ZN(new_n1203));
  NOR3_X1   g778(.A1(new_n1195), .A2(new_n1200), .A3(G1996), .ZN(new_n1204));
  XOR2_X1   g779(.A(new_n1204), .B(KEYINPUT126), .Z(new_n1205));
  OR3_X1    g780(.A1(new_n1202), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(KEYINPUT47), .ZN(new_n1207));
  OR2_X1    g782(.A1(new_n1206), .A2(KEYINPUT47), .ZN(new_n1208));
  AOI211_X1 g783(.A(new_n1194), .B(new_n1199), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g784(.A1(new_n1191), .A2(new_n1209), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g785(.A1(new_n649), .A2(new_n662), .ZN(new_n1212));
  AOI21_X1  g786(.A(new_n1212), .B1(new_n921), .B2(new_n922), .ZN(new_n1213));
  NAND4_X1  g787(.A1(new_n993), .A2(new_n460), .A3(new_n682), .A4(new_n1213), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n1214), .A2(KEYINPUT127), .ZN(new_n1215));
  INV_X1    g789(.A(new_n460), .ZN(new_n1216));
  AOI21_X1  g790(.A(new_n1216), .B1(new_n991), .B2(new_n992), .ZN(new_n1217));
  INV_X1    g791(.A(KEYINPUT127), .ZN(new_n1218));
  NAND4_X1  g792(.A1(new_n1217), .A2(new_n1218), .A3(new_n682), .A4(new_n1213), .ZN(new_n1219));
  AND2_X1   g793(.A1(new_n1215), .A2(new_n1219), .ZN(G308));
  NAND2_X1  g794(.A1(new_n1215), .A2(new_n1219), .ZN(G225));
endmodule


