

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U547 ( .A(KEYINPUT28), .ZN(n682) );
  NOR2_X1 U548 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U549 ( .A1(G651), .A2(n634), .ZN(n633) );
  AND2_X1 U550 ( .A1(G2104), .A2(G2105), .ZN(n881) );
  NAND2_X1 U551 ( .A1(n881), .A2(G113), .ZN(n522) );
  XNOR2_X1 U552 ( .A(KEYINPUT65), .B(KEYINPUT17), .ZN(n514) );
  NOR2_X1 U553 ( .A1(G2104), .A2(G2105), .ZN(n513) );
  XNOR2_X2 U554 ( .A(n514), .B(n513), .ZN(n877) );
  NAND2_X1 U555 ( .A1(G137), .A2(n877), .ZN(n516) );
  INV_X1 U556 ( .A(G2104), .ZN(n517) );
  AND2_X1 U557 ( .A1(n517), .A2(G2105), .ZN(n884) );
  NAND2_X1 U558 ( .A1(G125), .A2(n884), .ZN(n515) );
  NAND2_X1 U559 ( .A1(n516), .A2(n515), .ZN(n520) );
  NOR2_X4 U560 ( .A1(G2105), .A2(n517), .ZN(n876) );
  NAND2_X1 U561 ( .A1(G101), .A2(n876), .ZN(n518) );
  XNOR2_X1 U562 ( .A(KEYINPUT23), .B(n518), .ZN(n519) );
  NOR2_X1 U563 ( .A1(n520), .A2(n519), .ZN(n521) );
  NAND2_X1 U564 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X2 U565 ( .A(KEYINPUT64), .B(n523), .Z(G160) );
  XOR2_X1 U566 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  INV_X1 U567 ( .A(G651), .ZN(n532) );
  NOR2_X1 U568 ( .A1(n634), .A2(n532), .ZN(n625) );
  NAND2_X1 U569 ( .A1(G76), .A2(n625), .ZN(n528) );
  XOR2_X1 U570 ( .A(KEYINPUT4), .B(KEYINPUT75), .Z(n525) );
  NOR2_X1 U571 ( .A1(G651), .A2(G543), .ZN(n624) );
  NAND2_X1 U572 ( .A1(G89), .A2(n624), .ZN(n524) );
  XNOR2_X1 U573 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U574 ( .A(KEYINPUT74), .B(n526), .ZN(n527) );
  NAND2_X1 U575 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U576 ( .A(n529), .B(KEYINPUT76), .ZN(n530) );
  XNOR2_X1 U577 ( .A(KEYINPUT5), .B(n530), .ZN(n538) );
  NAND2_X1 U578 ( .A1(n633), .A2(G51), .ZN(n531) );
  XOR2_X1 U579 ( .A(KEYINPUT77), .B(n531), .Z(n535) );
  NOR2_X1 U580 ( .A1(G543), .A2(n532), .ZN(n533) );
  XOR2_X1 U581 ( .A(KEYINPUT1), .B(n533), .Z(n638) );
  NAND2_X1 U582 ( .A1(n638), .A2(G63), .ZN(n534) );
  NAND2_X1 U583 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U584 ( .A(KEYINPUT6), .B(n536), .Z(n537) );
  NAND2_X1 U585 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U586 ( .A(n539), .B(KEYINPUT7), .ZN(n540) );
  XNOR2_X1 U587 ( .A(KEYINPUT78), .B(n540), .ZN(G168) );
  XOR2_X1 U588 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U589 ( .A1(G85), .A2(n624), .ZN(n542) );
  NAND2_X1 U590 ( .A1(G72), .A2(n625), .ZN(n541) );
  NAND2_X1 U591 ( .A1(n542), .A2(n541), .ZN(n546) );
  NAND2_X1 U592 ( .A1(G60), .A2(n638), .ZN(n544) );
  NAND2_X1 U593 ( .A1(G47), .A2(n633), .ZN(n543) );
  NAND2_X1 U594 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U595 ( .A1(n546), .A2(n545), .ZN(G290) );
  NAND2_X1 U596 ( .A1(G52), .A2(n633), .ZN(n547) );
  XOR2_X1 U597 ( .A(KEYINPUT66), .B(n547), .Z(n554) );
  NAND2_X1 U598 ( .A1(G90), .A2(n624), .ZN(n549) );
  NAND2_X1 U599 ( .A1(G77), .A2(n625), .ZN(n548) );
  NAND2_X1 U600 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U601 ( .A(n550), .B(KEYINPUT9), .ZN(n552) );
  NAND2_X1 U602 ( .A1(G64), .A2(n638), .ZN(n551) );
  NAND2_X1 U603 ( .A1(n552), .A2(n551), .ZN(n553) );
  NOR2_X1 U604 ( .A1(n554), .A2(n553), .ZN(G171) );
  INV_X1 U605 ( .A(G57), .ZN(G237) );
  INV_X1 U606 ( .A(G108), .ZN(G238) );
  INV_X1 U607 ( .A(G120), .ZN(G236) );
  NAND2_X1 U608 ( .A1(G94), .A2(G452), .ZN(n555) );
  XNOR2_X1 U609 ( .A(n555), .B(KEYINPUT67), .ZN(G173) );
  NAND2_X1 U610 ( .A1(G7), .A2(G661), .ZN(n556) );
  XNOR2_X1 U611 ( .A(n556), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U612 ( .A(G223), .ZN(n813) );
  NAND2_X1 U613 ( .A1(n813), .A2(G567), .ZN(n557) );
  XOR2_X1 U614 ( .A(KEYINPUT11), .B(n557), .Z(G234) );
  XOR2_X1 U615 ( .A(G860), .B(KEYINPUT72), .Z(n590) );
  XOR2_X1 U616 ( .A(KEYINPUT70), .B(KEYINPUT14), .Z(n559) );
  NAND2_X1 U617 ( .A1(G56), .A2(n638), .ZN(n558) );
  XNOR2_X1 U618 ( .A(n559), .B(n558), .ZN(n566) );
  XNOR2_X1 U619 ( .A(KEYINPUT71), .B(KEYINPUT13), .ZN(n564) );
  NAND2_X1 U620 ( .A1(n624), .A2(G81), .ZN(n560) );
  XNOR2_X1 U621 ( .A(n560), .B(KEYINPUT12), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G68), .A2(n625), .ZN(n561) );
  NAND2_X1 U623 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U624 ( .A(n564), .B(n563), .ZN(n565) );
  NOR2_X1 U625 ( .A1(n566), .A2(n565), .ZN(n568) );
  NAND2_X1 U626 ( .A1(n633), .A2(G43), .ZN(n567) );
  NAND2_X1 U627 ( .A1(n568), .A2(n567), .ZN(n940) );
  OR2_X1 U628 ( .A1(n590), .A2(n940), .ZN(G153) );
  INV_X1 U629 ( .A(G171), .ZN(G301) );
  NAND2_X1 U630 ( .A1(G868), .A2(G301), .ZN(n578) );
  NAND2_X1 U631 ( .A1(G66), .A2(n638), .ZN(n570) );
  NAND2_X1 U632 ( .A1(G92), .A2(n624), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G79), .A2(n625), .ZN(n572) );
  NAND2_X1 U635 ( .A1(G54), .A2(n633), .ZN(n571) );
  NAND2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U637 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U638 ( .A(KEYINPUT15), .B(n575), .Z(n576) );
  XNOR2_X1 U639 ( .A(KEYINPUT73), .B(n576), .ZN(n933) );
  INV_X1 U640 ( .A(G868), .ZN(n650) );
  NAND2_X1 U641 ( .A1(n933), .A2(n650), .ZN(n577) );
  NAND2_X1 U642 ( .A1(n578), .A2(n577), .ZN(G284) );
  NAND2_X1 U643 ( .A1(n633), .A2(G53), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n579), .B(KEYINPUT68), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G65), .A2(n638), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(KEYINPUT69), .B(n582), .ZN(n586) );
  NAND2_X1 U648 ( .A1(G91), .A2(n624), .ZN(n584) );
  NAND2_X1 U649 ( .A1(G78), .A2(n625), .ZN(n583) );
  AND2_X1 U650 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(G299) );
  NOR2_X1 U652 ( .A1(G286), .A2(n650), .ZN(n587) );
  XOR2_X1 U653 ( .A(KEYINPUT79), .B(n587), .Z(n589) );
  NOR2_X1 U654 ( .A1(G868), .A2(G299), .ZN(n588) );
  NOR2_X1 U655 ( .A1(n589), .A2(n588), .ZN(G297) );
  NAND2_X1 U656 ( .A1(n590), .A2(G559), .ZN(n591) );
  INV_X1 U657 ( .A(n933), .ZN(n608) );
  NAND2_X1 U658 ( .A1(n591), .A2(n608), .ZN(n592) );
  XNOR2_X1 U659 ( .A(n592), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U660 ( .A1(G868), .A2(n940), .ZN(n593) );
  XNOR2_X1 U661 ( .A(KEYINPUT80), .B(n593), .ZN(n596) );
  NAND2_X1 U662 ( .A1(G868), .A2(n608), .ZN(n594) );
  NOR2_X1 U663 ( .A1(G559), .A2(n594), .ZN(n595) );
  NOR2_X1 U664 ( .A1(n596), .A2(n595), .ZN(G282) );
  XOR2_X1 U665 ( .A(KEYINPUT81), .B(KEYINPUT18), .Z(n598) );
  NAND2_X1 U666 ( .A1(G123), .A2(n884), .ZN(n597) );
  XNOR2_X1 U667 ( .A(n598), .B(n597), .ZN(n605) );
  NAND2_X1 U668 ( .A1(G99), .A2(n876), .ZN(n600) );
  NAND2_X1 U669 ( .A1(G135), .A2(n877), .ZN(n599) );
  NAND2_X1 U670 ( .A1(n600), .A2(n599), .ZN(n603) );
  NAND2_X1 U671 ( .A1(n881), .A2(G111), .ZN(n601) );
  XOR2_X1 U672 ( .A(KEYINPUT82), .B(n601), .Z(n602) );
  NOR2_X1 U673 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U674 ( .A1(n605), .A2(n604), .ZN(n993) );
  XNOR2_X1 U675 ( .A(G2096), .B(n993), .ZN(n606) );
  NOR2_X1 U676 ( .A1(n606), .A2(G2100), .ZN(n607) );
  XNOR2_X1 U677 ( .A(n607), .B(KEYINPUT83), .ZN(G156) );
  NAND2_X1 U678 ( .A1(G559), .A2(n608), .ZN(n609) );
  XNOR2_X1 U679 ( .A(n940), .B(n609), .ZN(n647) );
  NOR2_X1 U680 ( .A1(n647), .A2(G860), .ZN(n616) );
  NAND2_X1 U681 ( .A1(G67), .A2(n638), .ZN(n611) );
  NAND2_X1 U682 ( .A1(G93), .A2(n624), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U684 ( .A1(G80), .A2(n625), .ZN(n613) );
  NAND2_X1 U685 ( .A1(G55), .A2(n633), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  OR2_X1 U687 ( .A1(n615), .A2(n614), .ZN(n649) );
  XOR2_X1 U688 ( .A(n616), .B(n649), .Z(G145) );
  NAND2_X1 U689 ( .A1(G61), .A2(n638), .ZN(n618) );
  NAND2_X1 U690 ( .A1(G86), .A2(n624), .ZN(n617) );
  NAND2_X1 U691 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U692 ( .A1(n625), .A2(G73), .ZN(n619) );
  XOR2_X1 U693 ( .A(KEYINPUT2), .B(n619), .Z(n620) );
  NOR2_X1 U694 ( .A1(n621), .A2(n620), .ZN(n623) );
  NAND2_X1 U695 ( .A1(n633), .A2(G48), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n623), .A2(n622), .ZN(G305) );
  NAND2_X1 U697 ( .A1(G88), .A2(n624), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G75), .A2(n625), .ZN(n626) );
  NAND2_X1 U699 ( .A1(n627), .A2(n626), .ZN(n631) );
  NAND2_X1 U700 ( .A1(G62), .A2(n638), .ZN(n629) );
  NAND2_X1 U701 ( .A1(G50), .A2(n633), .ZN(n628) );
  NAND2_X1 U702 ( .A1(n629), .A2(n628), .ZN(n630) );
  NOR2_X1 U703 ( .A1(n631), .A2(n630), .ZN(G166) );
  NAND2_X1 U704 ( .A1(G74), .A2(G651), .ZN(n632) );
  XNOR2_X1 U705 ( .A(n632), .B(KEYINPUT84), .ZN(n640) );
  NAND2_X1 U706 ( .A1(G49), .A2(n633), .ZN(n636) );
  NAND2_X1 U707 ( .A1(G87), .A2(n634), .ZN(n635) );
  NAND2_X1 U708 ( .A1(n636), .A2(n635), .ZN(n637) );
  NOR2_X1 U709 ( .A1(n638), .A2(n637), .ZN(n639) );
  NAND2_X1 U710 ( .A1(n640), .A2(n639), .ZN(G288) );
  XOR2_X1 U711 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n642) );
  INV_X1 U712 ( .A(G299), .ZN(n685) );
  XNOR2_X1 U713 ( .A(n685), .B(G166), .ZN(n641) );
  XNOR2_X1 U714 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U715 ( .A(n649), .B(n643), .ZN(n644) );
  XNOR2_X1 U716 ( .A(G305), .B(n644), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n645), .B(G290), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n646), .B(G288), .ZN(n896) );
  XOR2_X1 U719 ( .A(n647), .B(n896), .Z(n648) );
  NAND2_X1 U720 ( .A1(n648), .A2(G868), .ZN(n652) );
  NAND2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U722 ( .A1(n652), .A2(n651), .ZN(G295) );
  NAND2_X1 U723 ( .A1(G2078), .A2(G2084), .ZN(n653) );
  XOR2_X1 U724 ( .A(KEYINPUT20), .B(n653), .Z(n654) );
  NAND2_X1 U725 ( .A1(G2090), .A2(n654), .ZN(n655) );
  XNOR2_X1 U726 ( .A(KEYINPUT21), .B(n655), .ZN(n656) );
  NAND2_X1 U727 ( .A1(n656), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U728 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U729 ( .A1(G236), .A2(G238), .ZN(n657) );
  NAND2_X1 U730 ( .A1(G69), .A2(n657), .ZN(n658) );
  NOR2_X1 U731 ( .A1(n658), .A2(G237), .ZN(n659) );
  XNOR2_X1 U732 ( .A(n659), .B(KEYINPUT89), .ZN(n818) );
  NAND2_X1 U733 ( .A1(n818), .A2(G567), .ZN(n667) );
  NAND2_X1 U734 ( .A1(G132), .A2(G82), .ZN(n660) );
  XNOR2_X1 U735 ( .A(n660), .B(KEYINPUT86), .ZN(n661) );
  XNOR2_X1 U736 ( .A(n661), .B(KEYINPUT22), .ZN(n662) );
  NOR2_X1 U737 ( .A1(G218), .A2(n662), .ZN(n663) );
  XOR2_X1 U738 ( .A(KEYINPUT87), .B(n663), .Z(n664) );
  NAND2_X1 U739 ( .A1(n664), .A2(G96), .ZN(n665) );
  XNOR2_X1 U740 ( .A(n665), .B(KEYINPUT88), .ZN(n819) );
  NAND2_X1 U741 ( .A1(n819), .A2(G2106), .ZN(n666) );
  NAND2_X1 U742 ( .A1(n667), .A2(n666), .ZN(n820) );
  NAND2_X1 U743 ( .A1(G483), .A2(G661), .ZN(n668) );
  NOR2_X1 U744 ( .A1(n820), .A2(n668), .ZN(n817) );
  NAND2_X1 U745 ( .A1(n817), .A2(G36), .ZN(G176) );
  NAND2_X1 U746 ( .A1(n876), .A2(G102), .ZN(n669) );
  XNOR2_X1 U747 ( .A(n669), .B(KEYINPUT90), .ZN(n671) );
  NAND2_X1 U748 ( .A1(G138), .A2(n877), .ZN(n670) );
  NAND2_X1 U749 ( .A1(n671), .A2(n670), .ZN(n675) );
  NAND2_X1 U750 ( .A1(G126), .A2(n884), .ZN(n673) );
  NAND2_X1 U751 ( .A1(G114), .A2(n881), .ZN(n672) );
  NAND2_X1 U752 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U753 ( .A1(n675), .A2(n674), .ZN(G164) );
  XNOR2_X1 U754 ( .A(KEYINPUT91), .B(G166), .ZN(G303) );
  NOR2_X1 U755 ( .A1(G164), .A2(G1384), .ZN(n763) );
  AND2_X1 U756 ( .A1(G40), .A2(n763), .ZN(n676) );
  NAND2_X2 U757 ( .A1(G160), .A2(n676), .ZN(n720) );
  NAND2_X1 U758 ( .A1(G1956), .A2(n720), .ZN(n680) );
  INV_X1 U759 ( .A(n720), .ZN(n677) );
  NAND2_X1 U760 ( .A1(n677), .A2(G2072), .ZN(n678) );
  XOR2_X1 U761 ( .A(n678), .B(KEYINPUT27), .Z(n679) );
  NAND2_X1 U762 ( .A1(n680), .A2(n679), .ZN(n681) );
  XOR2_X1 U763 ( .A(n681), .B(KEYINPUT98), .Z(n684) );
  NOR2_X1 U764 ( .A1(n685), .A2(n684), .ZN(n683) );
  XNOR2_X1 U765 ( .A(n683), .B(n682), .ZN(n700) );
  NAND2_X1 U766 ( .A1(n685), .A2(n684), .ZN(n698) );
  INV_X1 U767 ( .A(n720), .ZN(n703) );
  AND2_X1 U768 ( .A1(n703), .A2(G1996), .ZN(n686) );
  XOR2_X1 U769 ( .A(n686), .B(KEYINPUT26), .Z(n688) );
  NAND2_X1 U770 ( .A1(n720), .A2(G1341), .ZN(n687) );
  NAND2_X1 U771 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U772 ( .A1(n940), .A2(n689), .ZN(n693) );
  NAND2_X1 U773 ( .A1(G1348), .A2(n720), .ZN(n691) );
  NAND2_X1 U774 ( .A1(G2067), .A2(n703), .ZN(n690) );
  NAND2_X1 U775 ( .A1(n691), .A2(n690), .ZN(n694) );
  NOR2_X1 U776 ( .A1(n933), .A2(n694), .ZN(n692) );
  OR2_X1 U777 ( .A1(n693), .A2(n692), .ZN(n696) );
  NAND2_X1 U778 ( .A1(n933), .A2(n694), .ZN(n695) );
  NAND2_X1 U779 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U780 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U781 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U782 ( .A(n701), .B(KEYINPUT29), .ZN(n708) );
  XNOR2_X1 U783 ( .A(G2078), .B(KEYINPUT96), .ZN(n702) );
  XNOR2_X1 U784 ( .A(n702), .B(KEYINPUT25), .ZN(n914) );
  NOR2_X1 U785 ( .A1(n914), .A2(n720), .ZN(n705) );
  INV_X1 U786 ( .A(G1961), .ZN(n964) );
  NOR2_X1 U787 ( .A1(n703), .A2(n964), .ZN(n704) );
  NOR2_X1 U788 ( .A1(n705), .A2(n704), .ZN(n713) );
  AND2_X1 U789 ( .A1(G171), .A2(n713), .ZN(n706) );
  XOR2_X1 U790 ( .A(KEYINPUT97), .B(n706), .Z(n707) );
  XNOR2_X1 U791 ( .A(n709), .B(KEYINPUT99), .ZN(n718) );
  NAND2_X1 U792 ( .A1(G8), .A2(n720), .ZN(n754) );
  NOR2_X1 U793 ( .A1(G1966), .A2(n754), .ZN(n732) );
  NOR2_X1 U794 ( .A1(G2084), .A2(n720), .ZN(n729) );
  NOR2_X1 U795 ( .A1(n732), .A2(n729), .ZN(n710) );
  NAND2_X1 U796 ( .A1(G8), .A2(n710), .ZN(n711) );
  XNOR2_X1 U797 ( .A(KEYINPUT30), .B(n711), .ZN(n712) );
  NOR2_X1 U798 ( .A1(G168), .A2(n712), .ZN(n715) );
  NOR2_X1 U799 ( .A1(G171), .A2(n713), .ZN(n714) );
  NOR2_X1 U800 ( .A1(n715), .A2(n714), .ZN(n716) );
  XOR2_X1 U801 ( .A(KEYINPUT31), .B(n716), .Z(n717) );
  NAND2_X1 U802 ( .A1(n718), .A2(n717), .ZN(n730) );
  NAND2_X1 U803 ( .A1(n730), .A2(G286), .ZN(n719) );
  XNOR2_X1 U804 ( .A(n719), .B(KEYINPUT100), .ZN(n725) );
  NOR2_X1 U805 ( .A1(G1971), .A2(n754), .ZN(n722) );
  NOR2_X1 U806 ( .A1(G2090), .A2(n720), .ZN(n721) );
  NOR2_X1 U807 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U808 ( .A1(n723), .A2(G303), .ZN(n724) );
  NAND2_X1 U809 ( .A1(n725), .A2(n724), .ZN(n726) );
  NAND2_X1 U810 ( .A1(n726), .A2(G8), .ZN(n728) );
  XOR2_X1 U811 ( .A(KEYINPUT32), .B(KEYINPUT101), .Z(n727) );
  XNOR2_X1 U812 ( .A(n728), .B(n727), .ZN(n746) );
  NAND2_X1 U813 ( .A1(G8), .A2(n729), .ZN(n734) );
  INV_X1 U814 ( .A(n730), .ZN(n731) );
  NOR2_X1 U815 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U816 ( .A1(n734), .A2(n733), .ZN(n744) );
  NAND2_X1 U817 ( .A1(n746), .A2(n744), .ZN(n737) );
  NOR2_X1 U818 ( .A1(G2090), .A2(G303), .ZN(n735) );
  NAND2_X1 U819 ( .A1(G8), .A2(n735), .ZN(n736) );
  NAND2_X1 U820 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U821 ( .A1(n738), .A2(n754), .ZN(n743) );
  NOR2_X1 U822 ( .A1(G1981), .A2(G305), .ZN(n739) );
  XNOR2_X1 U823 ( .A(n739), .B(KEYINPUT24), .ZN(n740) );
  XNOR2_X1 U824 ( .A(n740), .B(KEYINPUT95), .ZN(n741) );
  OR2_X1 U825 ( .A1(n741), .A2(n754), .ZN(n742) );
  AND2_X1 U826 ( .A1(n743), .A2(n742), .ZN(n761) );
  NAND2_X1 U827 ( .A1(G1976), .A2(G288), .ZN(n747) );
  AND2_X1 U828 ( .A1(n744), .A2(n747), .ZN(n745) );
  NAND2_X1 U829 ( .A1(n746), .A2(n745), .ZN(n752) );
  INV_X1 U830 ( .A(n747), .ZN(n930) );
  NOR2_X1 U831 ( .A1(G1976), .A2(G288), .ZN(n753) );
  NOR2_X1 U832 ( .A1(G1971), .A2(G303), .ZN(n748) );
  NOR2_X1 U833 ( .A1(n753), .A2(n748), .ZN(n937) );
  OR2_X1 U834 ( .A1(n930), .A2(n937), .ZN(n749) );
  NOR2_X1 U835 ( .A1(n754), .A2(n749), .ZN(n750) );
  NOR2_X1 U836 ( .A1(n750), .A2(KEYINPUT33), .ZN(n751) );
  NAND2_X1 U837 ( .A1(n752), .A2(n751), .ZN(n759) );
  NAND2_X1 U838 ( .A1(n753), .A2(KEYINPUT33), .ZN(n755) );
  NOR2_X1 U839 ( .A1(n755), .A2(n754), .ZN(n757) );
  XOR2_X1 U840 ( .A(G1981), .B(G305), .Z(n943) );
  INV_X1 U841 ( .A(n943), .ZN(n756) );
  NOR2_X1 U842 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U843 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U844 ( .A1(n761), .A2(n760), .ZN(n794) );
  NAND2_X1 U845 ( .A1(G40), .A2(G160), .ZN(n762) );
  NOR2_X1 U846 ( .A1(n763), .A2(n762), .ZN(n809) );
  NAND2_X1 U847 ( .A1(G128), .A2(n884), .ZN(n765) );
  NAND2_X1 U848 ( .A1(G116), .A2(n881), .ZN(n764) );
  NAND2_X1 U849 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U850 ( .A(n766), .B(KEYINPUT35), .ZN(n771) );
  NAND2_X1 U851 ( .A1(G104), .A2(n876), .ZN(n768) );
  NAND2_X1 U852 ( .A1(G140), .A2(n877), .ZN(n767) );
  NAND2_X1 U853 ( .A1(n768), .A2(n767), .ZN(n769) );
  XOR2_X1 U854 ( .A(KEYINPUT34), .B(n769), .Z(n770) );
  NAND2_X1 U855 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U856 ( .A(n772), .B(KEYINPUT36), .ZN(n890) );
  XOR2_X1 U857 ( .A(KEYINPUT37), .B(G2067), .Z(n805) );
  NAND2_X1 U858 ( .A1(n890), .A2(n805), .ZN(n773) );
  XOR2_X1 U859 ( .A(KEYINPUT92), .B(n773), .Z(n1000) );
  NAND2_X1 U860 ( .A1(n809), .A2(n1000), .ZN(n803) );
  INV_X1 U861 ( .A(n803), .ZN(n792) );
  XNOR2_X1 U862 ( .A(KEYINPUT94), .B(n809), .ZN(n789) );
  NAND2_X1 U863 ( .A1(G129), .A2(n884), .ZN(n775) );
  NAND2_X1 U864 ( .A1(G141), .A2(n877), .ZN(n774) );
  NAND2_X1 U865 ( .A1(n775), .A2(n774), .ZN(n778) );
  NAND2_X1 U866 ( .A1(n876), .A2(G105), .ZN(n776) );
  XOR2_X1 U867 ( .A(KEYINPUT38), .B(n776), .Z(n777) );
  NOR2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n881), .A2(G117), .ZN(n779) );
  NAND2_X1 U870 ( .A1(n780), .A2(n779), .ZN(n889) );
  NAND2_X1 U871 ( .A1(G1996), .A2(n889), .ZN(n788) );
  XNOR2_X1 U872 ( .A(KEYINPUT93), .B(G1991), .ZN(n915) );
  NAND2_X1 U873 ( .A1(G95), .A2(n876), .ZN(n782) );
  NAND2_X1 U874 ( .A1(G119), .A2(n884), .ZN(n781) );
  NAND2_X1 U875 ( .A1(n782), .A2(n781), .ZN(n786) );
  NAND2_X1 U876 ( .A1(G131), .A2(n877), .ZN(n784) );
  NAND2_X1 U877 ( .A1(G107), .A2(n881), .ZN(n783) );
  NAND2_X1 U878 ( .A1(n784), .A2(n783), .ZN(n785) );
  NOR2_X1 U879 ( .A1(n786), .A2(n785), .ZN(n862) );
  OR2_X1 U880 ( .A1(n915), .A2(n862), .ZN(n787) );
  NAND2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n996) );
  NAND2_X1 U882 ( .A1(n789), .A2(n996), .ZN(n798) );
  XNOR2_X1 U883 ( .A(G1986), .B(G290), .ZN(n929) );
  NAND2_X1 U884 ( .A1(n809), .A2(n929), .ZN(n790) );
  NAND2_X1 U885 ( .A1(n798), .A2(n790), .ZN(n791) );
  NOR2_X1 U886 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U887 ( .A1(n794), .A2(n793), .ZN(n795) );
  XNOR2_X1 U888 ( .A(n795), .B(KEYINPUT102), .ZN(n811) );
  NOR2_X1 U889 ( .A1(G1996), .A2(n889), .ZN(n984) );
  NOR2_X1 U890 ( .A1(G1986), .A2(G290), .ZN(n796) );
  XNOR2_X1 U891 ( .A(KEYINPUT103), .B(n796), .ZN(n797) );
  NAND2_X1 U892 ( .A1(n862), .A2(n915), .ZN(n994) );
  NAND2_X1 U893 ( .A1(n797), .A2(n994), .ZN(n799) );
  NAND2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U895 ( .A(KEYINPUT104), .B(n800), .Z(n801) );
  NOR2_X1 U896 ( .A1(n984), .A2(n801), .ZN(n802) );
  XNOR2_X1 U897 ( .A(n802), .B(KEYINPUT39), .ZN(n804) );
  NAND2_X1 U898 ( .A1(n804), .A2(n803), .ZN(n807) );
  NOR2_X1 U899 ( .A1(n805), .A2(n890), .ZN(n806) );
  XNOR2_X1 U900 ( .A(n806), .B(KEYINPUT105), .ZN(n1003) );
  NAND2_X1 U901 ( .A1(n807), .A2(n1003), .ZN(n808) );
  NAND2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n810) );
  NAND2_X1 U903 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U904 ( .A(n812), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U905 ( .A1(G2106), .A2(n813), .ZN(G217) );
  NAND2_X1 U906 ( .A1(G15), .A2(G2), .ZN(n814) );
  XOR2_X1 U907 ( .A(KEYINPUT108), .B(n814), .Z(n815) );
  NAND2_X1 U908 ( .A1(G661), .A2(n815), .ZN(G259) );
  NAND2_X1 U909 ( .A1(G3), .A2(G1), .ZN(n816) );
  NAND2_X1 U910 ( .A1(n817), .A2(n816), .ZN(G188) );
  XNOR2_X1 U911 ( .A(G96), .B(KEYINPUT109), .ZN(G221) );
  INV_X1 U913 ( .A(G132), .ZN(G219) );
  INV_X1 U914 ( .A(G82), .ZN(G220) );
  NOR2_X1 U915 ( .A1(n819), .A2(n818), .ZN(G325) );
  INV_X1 U916 ( .A(G325), .ZN(G261) );
  INV_X1 U917 ( .A(n820), .ZN(G319) );
  XNOR2_X1 U918 ( .A(G2454), .B(G2435), .ZN(n829) );
  XNOR2_X1 U919 ( .A(KEYINPUT106), .B(G2427), .ZN(n827) );
  XOR2_X1 U920 ( .A(G2430), .B(G2446), .Z(n822) );
  XNOR2_X1 U921 ( .A(G2443), .B(G2451), .ZN(n821) );
  XNOR2_X1 U922 ( .A(n822), .B(n821), .ZN(n823) );
  XOR2_X1 U923 ( .A(n823), .B(G2438), .Z(n825) );
  XNOR2_X1 U924 ( .A(G1341), .B(G1348), .ZN(n824) );
  XNOR2_X1 U925 ( .A(n825), .B(n824), .ZN(n826) );
  XNOR2_X1 U926 ( .A(n827), .B(n826), .ZN(n828) );
  XNOR2_X1 U927 ( .A(n829), .B(n828), .ZN(n830) );
  NAND2_X1 U928 ( .A1(n830), .A2(G14), .ZN(n831) );
  XNOR2_X1 U929 ( .A(KEYINPUT107), .B(n831), .ZN(G401) );
  XNOR2_X1 U930 ( .A(G1961), .B(KEYINPUT41), .ZN(n841) );
  XOR2_X1 U931 ( .A(G1976), .B(G1971), .Z(n833) );
  XNOR2_X1 U932 ( .A(G1986), .B(G1956), .ZN(n832) );
  XNOR2_X1 U933 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U934 ( .A(G1981), .B(G1966), .Z(n835) );
  XNOR2_X1 U935 ( .A(G1996), .B(G1991), .ZN(n834) );
  XNOR2_X1 U936 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U937 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U938 ( .A(KEYINPUT112), .B(G2474), .ZN(n838) );
  XNOR2_X1 U939 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(G229) );
  XOR2_X1 U941 ( .A(KEYINPUT43), .B(KEYINPUT111), .Z(n843) );
  XNOR2_X1 U942 ( .A(KEYINPUT110), .B(G2678), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U944 ( .A(KEYINPUT42), .B(G2090), .Z(n845) );
  XNOR2_X1 U945 ( .A(G2067), .B(G2072), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U947 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U948 ( .A(G2096), .B(G2100), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n851) );
  XOR2_X1 U950 ( .A(G2078), .B(G2084), .Z(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(G227) );
  NAND2_X1 U952 ( .A1(n877), .A2(G136), .ZN(n852) );
  XNOR2_X1 U953 ( .A(KEYINPUT113), .B(n852), .ZN(n855) );
  NAND2_X1 U954 ( .A1(n884), .A2(G124), .ZN(n853) );
  XOR2_X1 U955 ( .A(KEYINPUT44), .B(n853), .Z(n854) );
  NOR2_X1 U956 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n856), .B(KEYINPUT114), .ZN(n858) );
  NAND2_X1 U958 ( .A1(G112), .A2(n881), .ZN(n857) );
  NAND2_X1 U959 ( .A1(n858), .A2(n857), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G100), .A2(n876), .ZN(n859) );
  XNOR2_X1 U961 ( .A(KEYINPUT115), .B(n859), .ZN(n860) );
  NOR2_X1 U962 ( .A1(n861), .A2(n860), .ZN(G162) );
  XNOR2_X1 U963 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n864) );
  XNOR2_X1 U964 ( .A(G160), .B(n862), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U966 ( .A(n993), .B(n865), .ZN(n875) );
  NAND2_X1 U967 ( .A1(G127), .A2(n884), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G115), .A2(n881), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U970 ( .A(n868), .B(KEYINPUT47), .ZN(n870) );
  NAND2_X1 U971 ( .A1(G103), .A2(n876), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n873) );
  NAND2_X1 U973 ( .A1(G139), .A2(n877), .ZN(n871) );
  XNOR2_X1 U974 ( .A(KEYINPUT117), .B(n871), .ZN(n872) );
  NOR2_X1 U975 ( .A1(n873), .A2(n872), .ZN(n987) );
  XNOR2_X1 U976 ( .A(G162), .B(n987), .ZN(n874) );
  XNOR2_X1 U977 ( .A(n875), .B(n874), .ZN(n894) );
  NAND2_X1 U978 ( .A1(G106), .A2(n876), .ZN(n879) );
  NAND2_X1 U979 ( .A1(G142), .A2(n877), .ZN(n878) );
  NAND2_X1 U980 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n880), .B(KEYINPUT45), .ZN(n883) );
  NAND2_X1 U982 ( .A1(G118), .A2(n881), .ZN(n882) );
  NAND2_X1 U983 ( .A1(n883), .A2(n882), .ZN(n887) );
  NAND2_X1 U984 ( .A1(n884), .A2(G130), .ZN(n885) );
  XOR2_X1 U985 ( .A(KEYINPUT116), .B(n885), .Z(n886) );
  NOR2_X1 U986 ( .A1(n887), .A2(n886), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n889), .B(n888), .ZN(n892) );
  XNOR2_X1 U988 ( .A(G164), .B(n890), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U990 ( .A(n894), .B(n893), .Z(n895) );
  NOR2_X1 U991 ( .A1(G37), .A2(n895), .ZN(G395) );
  XNOR2_X1 U992 ( .A(KEYINPUT118), .B(n933), .ZN(n899) );
  XNOR2_X1 U993 ( .A(G171), .B(n896), .ZN(n897) );
  XNOR2_X1 U994 ( .A(n897), .B(n940), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U996 ( .A(n900), .B(G286), .Z(n901) );
  NOR2_X1 U997 ( .A1(G37), .A2(n901), .ZN(G397) );
  NOR2_X1 U998 ( .A1(G229), .A2(G227), .ZN(n902) );
  XOR2_X1 U999 ( .A(KEYINPUT49), .B(n902), .Z(n903) );
  XNOR2_X1 U1000 ( .A(n903), .B(KEYINPUT119), .ZN(n904) );
  NOR2_X1 U1001 ( .A1(G401), .A2(n904), .ZN(n905) );
  AND2_X1 U1002 ( .A1(G319), .A2(n905), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(n907), .A2(n906), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  INV_X1 U1006 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1007 ( .A(KEYINPUT55), .B(KEYINPUT122), .Z(n1007) );
  XNOR2_X1 U1008 ( .A(G1996), .B(G32), .ZN(n909) );
  XNOR2_X1 U1009 ( .A(G33), .B(G2072), .ZN(n908) );
  NOR2_X1 U1010 ( .A1(n909), .A2(n908), .ZN(n910) );
  NAND2_X1 U1011 ( .A1(G28), .A2(n910), .ZN(n913) );
  XOR2_X1 U1012 ( .A(KEYINPUT123), .B(G2067), .Z(n911) );
  XNOR2_X1 U1013 ( .A(G26), .B(n911), .ZN(n912) );
  NOR2_X1 U1014 ( .A1(n913), .A2(n912), .ZN(n919) );
  XOR2_X1 U1015 ( .A(n914), .B(G27), .Z(n917) );
  XOR2_X1 U1016 ( .A(G25), .B(n915), .Z(n916) );
  NOR2_X1 U1017 ( .A1(n917), .A2(n916), .ZN(n918) );
  NAND2_X1 U1018 ( .A1(n919), .A2(n918), .ZN(n920) );
  XNOR2_X1 U1019 ( .A(n920), .B(KEYINPUT53), .ZN(n923) );
  XOR2_X1 U1020 ( .A(G2084), .B(G34), .Z(n921) );
  XNOR2_X1 U1021 ( .A(KEYINPUT54), .B(n921), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n923), .A2(n922), .ZN(n925) );
  XNOR2_X1 U1023 ( .A(G35), .B(G2090), .ZN(n924) );
  NOR2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(n1007), .B(n926), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(KEYINPUT124), .B(G29), .ZN(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n980) );
  XNOR2_X1 U1028 ( .A(G16), .B(KEYINPUT56), .ZN(n951) );
  NOR2_X1 U1029 ( .A1(n930), .A2(n929), .ZN(n932) );
  NAND2_X1 U1030 ( .A1(G1971), .A2(G303), .ZN(n931) );
  NAND2_X1 U1031 ( .A1(n932), .A2(n931), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(G1348), .B(n933), .ZN(n934) );
  NOR2_X1 U1033 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n939) );
  XNOR2_X1 U1035 ( .A(G1956), .B(G299), .ZN(n938) );
  NOR2_X1 U1036 ( .A1(n939), .A2(n938), .ZN(n949) );
  XOR2_X1 U1037 ( .A(n940), .B(G1341), .Z(n942) );
  XNOR2_X1 U1038 ( .A(G171), .B(G1961), .ZN(n941) );
  NAND2_X1 U1039 ( .A1(n942), .A2(n941), .ZN(n947) );
  XNOR2_X1 U1040 ( .A(G1966), .B(G168), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1042 ( .A(KEYINPUT57), .B(n945), .Z(n946) );
  NOR2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  NAND2_X1 U1044 ( .A1(n949), .A2(n948), .ZN(n950) );
  NAND2_X1 U1045 ( .A1(n951), .A2(n950), .ZN(n978) );
  INV_X1 U1046 ( .A(G16), .ZN(n976) );
  XNOR2_X1 U1047 ( .A(G1348), .B(KEYINPUT59), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(n952), .B(G4), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(G1341), .B(G19), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G1956), .B(G20), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n959) );
  XOR2_X1 U1053 ( .A(KEYINPUT125), .B(G1981), .Z(n957) );
  XNOR2_X1 U1054 ( .A(G6), .B(n957), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XOR2_X1 U1056 ( .A(KEYINPUT60), .B(n960), .Z(n962) );
  XNOR2_X1 U1057 ( .A(G1966), .B(G21), .ZN(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1059 ( .A(KEYINPUT126), .B(n963), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n964), .B(G5), .ZN(n965) );
  NAND2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n973) );
  XNOR2_X1 U1062 ( .A(G1971), .B(G22), .ZN(n968) );
  XNOR2_X1 U1063 ( .A(G23), .B(G1976), .ZN(n967) );
  NOR2_X1 U1064 ( .A1(n968), .A2(n967), .ZN(n970) );
  XOR2_X1 U1065 ( .A(G1986), .B(G24), .Z(n969) );
  NAND2_X1 U1066 ( .A1(n970), .A2(n969), .ZN(n971) );
  XNOR2_X1 U1067 ( .A(KEYINPUT58), .B(n971), .ZN(n972) );
  NOR2_X1 U1068 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(KEYINPUT61), .B(n974), .ZN(n975) );
  NAND2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n979) );
  NOR2_X1 U1072 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1073 ( .A1(G11), .A2(n981), .ZN(n982) );
  XNOR2_X1 U1074 ( .A(n982), .B(KEYINPUT127), .ZN(n1011) );
  XOR2_X1 U1075 ( .A(G2090), .B(G162), .Z(n983) );
  NOR2_X1 U1076 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1077 ( .A(KEYINPUT51), .B(n985), .Z(n986) );
  XOR2_X1 U1078 ( .A(KEYINPUT121), .B(n986), .Z(n992) );
  XOR2_X1 U1079 ( .A(G2072), .B(n987), .Z(n989) );
  XOR2_X1 U1080 ( .A(G164), .B(G2078), .Z(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1082 ( .A(KEYINPUT50), .B(n990), .ZN(n991) );
  NAND2_X1 U1083 ( .A1(n992), .A2(n991), .ZN(n1005) );
  XNOR2_X1 U1084 ( .A(G2084), .B(G160), .ZN(n998) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NOR2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1088 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1089 ( .A(n1001), .B(KEYINPUT120), .ZN(n1002) );
  NAND2_X1 U1090 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NOR2_X1 U1091 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1092 ( .A(KEYINPUT52), .B(n1006), .ZN(n1008) );
  NAND2_X1 U1093 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1094 ( .A1(n1009), .A2(G29), .ZN(n1010) );
  NAND2_X1 U1095 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1096 ( .A(KEYINPUT62), .B(n1012), .Z(G311) );
  INV_X1 U1097 ( .A(G311), .ZN(G150) );
endmodule

