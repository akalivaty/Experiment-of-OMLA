

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U558 ( .A(n531), .B(KEYINPUT65), .ZN(n999) );
  XNOR2_X1 U559 ( .A(n534), .B(n533), .ZN(n535) );
  INV_X1 U560 ( .A(KEYINPUT23), .ZN(n533) );
  NOR2_X1 U561 ( .A1(n739), .A2(n889), .ZN(n714) );
  NOR2_X1 U562 ( .A1(n779), .A2(n778), .ZN(n780) );
  INV_X1 U563 ( .A(G2104), .ZN(n532) );
  NOR2_X1 U564 ( .A1(G651), .A2(n622), .ZN(n645) );
  NOR2_X2 U565 ( .A1(G2105), .A2(n532), .ZN(n1004) );
  XNOR2_X1 U566 ( .A(KEYINPUT67), .B(KEYINPUT17), .ZN(n526) );
  NOR2_X1 U567 ( .A1(G2104), .A2(G2105), .ZN(n525) );
  XNOR2_X1 U568 ( .A(n526), .B(n525), .ZN(n527) );
  XNOR2_X1 U569 ( .A(KEYINPUT66), .B(n527), .ZN(n604) );
  NAND2_X1 U570 ( .A1(G137), .A2(n604), .ZN(n529) );
  AND2_X1 U571 ( .A1(G2104), .A2(G2105), .ZN(n998) );
  NAND2_X1 U572 ( .A1(n998), .A2(G113), .ZN(n528) );
  NAND2_X1 U573 ( .A1(n529), .A2(n528), .ZN(n530) );
  XNOR2_X1 U574 ( .A(KEYINPUT68), .B(n530), .ZN(n538) );
  NAND2_X1 U575 ( .A1(n532), .A2(G2105), .ZN(n531) );
  NAND2_X1 U576 ( .A1(n999), .A2(G125), .ZN(n536) );
  NAND2_X1 U577 ( .A1(G101), .A2(n1004), .ZN(n534) );
  NAND2_X1 U578 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U579 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X2 U580 ( .A(KEYINPUT64), .B(n539), .ZN(G160) );
  XNOR2_X1 U581 ( .A(G543), .B(KEYINPUT0), .ZN(n540) );
  XNOR2_X1 U582 ( .A(n540), .B(KEYINPUT69), .ZN(n622) );
  NAND2_X1 U583 ( .A1(G52), .A2(n645), .ZN(n543) );
  INV_X1 U584 ( .A(G651), .ZN(n544) );
  NOR2_X1 U585 ( .A1(G543), .A2(n544), .ZN(n541) );
  XOR2_X1 U586 ( .A(KEYINPUT1), .B(n541), .Z(n648) );
  NAND2_X1 U587 ( .A1(G64), .A2(n648), .ZN(n542) );
  NAND2_X1 U588 ( .A1(n543), .A2(n542), .ZN(n550) );
  NOR2_X1 U589 ( .A1(n622), .A2(n544), .ZN(n651) );
  NAND2_X1 U590 ( .A1(G77), .A2(n651), .ZN(n546) );
  NOR2_X1 U591 ( .A1(G651), .A2(G543), .ZN(n647) );
  NAND2_X1 U592 ( .A1(G90), .A2(n647), .ZN(n545) );
  NAND2_X1 U593 ( .A1(n546), .A2(n545), .ZN(n547) );
  XOR2_X1 U594 ( .A(KEYINPUT72), .B(n547), .Z(n548) );
  XNOR2_X1 U595 ( .A(KEYINPUT9), .B(n548), .ZN(n549) );
  NOR2_X1 U596 ( .A1(n550), .A2(n549), .ZN(G171) );
  AND2_X1 U597 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U598 ( .A(G120), .ZN(G236) );
  NAND2_X1 U599 ( .A1(n647), .A2(G89), .ZN(n551) );
  XNOR2_X1 U600 ( .A(n551), .B(KEYINPUT4), .ZN(n553) );
  NAND2_X1 U601 ( .A1(G76), .A2(n651), .ZN(n552) );
  NAND2_X1 U602 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U603 ( .A(n554), .B(KEYINPUT5), .ZN(n560) );
  XNOR2_X1 U604 ( .A(KEYINPUT6), .B(KEYINPUT79), .ZN(n558) );
  NAND2_X1 U605 ( .A1(G51), .A2(n645), .ZN(n556) );
  NAND2_X1 U606 ( .A1(G63), .A2(n648), .ZN(n555) );
  NAND2_X1 U607 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U608 ( .A(n558), .B(n557), .ZN(n559) );
  NAND2_X1 U609 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U610 ( .A(KEYINPUT7), .B(n561), .ZN(G168) );
  XOR2_X1 U611 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U612 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U613 ( .A(n562), .B(KEYINPUT76), .ZN(n563) );
  XNOR2_X1 U614 ( .A(KEYINPUT10), .B(n563), .ZN(G223) );
  INV_X1 U615 ( .A(G223), .ZN(n835) );
  NAND2_X1 U616 ( .A1(n835), .A2(G567), .ZN(n564) );
  XOR2_X1 U617 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  NAND2_X1 U618 ( .A1(G56), .A2(n648), .ZN(n565) );
  XOR2_X1 U619 ( .A(KEYINPUT14), .B(n565), .Z(n572) );
  NAND2_X1 U620 ( .A1(G81), .A2(n647), .ZN(n566) );
  XOR2_X1 U621 ( .A(KEYINPUT12), .B(n566), .Z(n567) );
  XNOR2_X1 U622 ( .A(n567), .B(KEYINPUT77), .ZN(n569) );
  NAND2_X1 U623 ( .A1(G68), .A2(n651), .ZN(n568) );
  NAND2_X1 U624 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U625 ( .A(KEYINPUT13), .B(n570), .Z(n571) );
  NOR2_X1 U626 ( .A1(n572), .A2(n571), .ZN(n574) );
  NAND2_X1 U627 ( .A1(n645), .A2(G43), .ZN(n573) );
  NAND2_X1 U628 ( .A1(n574), .A2(n573), .ZN(n1020) );
  INV_X1 U629 ( .A(G860), .ZN(n595) );
  OR2_X1 U630 ( .A1(n1020), .A2(n595), .ZN(G153) );
  INV_X1 U631 ( .A(G171), .ZN(G301) );
  NAND2_X1 U632 ( .A1(G92), .A2(n647), .ZN(n576) );
  NAND2_X1 U633 ( .A1(G66), .A2(n648), .ZN(n575) );
  NAND2_X1 U634 ( .A1(n576), .A2(n575), .ZN(n580) );
  NAND2_X1 U635 ( .A1(G79), .A2(n651), .ZN(n578) );
  NAND2_X1 U636 ( .A1(G54), .A2(n645), .ZN(n577) );
  NAND2_X1 U637 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U638 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U639 ( .A(KEYINPUT15), .B(n581), .Z(n582) );
  XNOR2_X1 U640 ( .A(KEYINPUT78), .B(n582), .ZN(n907) );
  INV_X1 U641 ( .A(n907), .ZN(n1017) );
  NOR2_X1 U642 ( .A1(n1017), .A2(G868), .ZN(n584) );
  INV_X1 U643 ( .A(G868), .ZN(n668) );
  NOR2_X1 U644 ( .A1(n668), .A2(G301), .ZN(n583) );
  NOR2_X1 U645 ( .A1(n584), .A2(n583), .ZN(G284) );
  NAND2_X1 U646 ( .A1(G65), .A2(n648), .ZN(n591) );
  NAND2_X1 U647 ( .A1(G78), .A2(n651), .ZN(n586) );
  NAND2_X1 U648 ( .A1(G53), .A2(n645), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U650 ( .A1(G91), .A2(n647), .ZN(n587) );
  XNOR2_X1 U651 ( .A(KEYINPUT73), .B(n587), .ZN(n588) );
  NOR2_X1 U652 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U653 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U654 ( .A(n592), .B(KEYINPUT74), .ZN(G299) );
  NOR2_X1 U655 ( .A1(G286), .A2(n668), .ZN(n594) );
  NOR2_X1 U656 ( .A1(G299), .A2(G868), .ZN(n593) );
  NOR2_X1 U657 ( .A1(n594), .A2(n593), .ZN(G297) );
  NAND2_X1 U658 ( .A1(n595), .A2(G559), .ZN(n596) );
  NAND2_X1 U659 ( .A1(n596), .A2(n907), .ZN(n597) );
  XNOR2_X1 U660 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U661 ( .A1(G868), .A2(n1020), .ZN(n600) );
  NAND2_X1 U662 ( .A1(n907), .A2(G868), .ZN(n598) );
  NOR2_X1 U663 ( .A1(G559), .A2(n598), .ZN(n599) );
  NOR2_X1 U664 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U665 ( .A1(G99), .A2(n1004), .ZN(n602) );
  NAND2_X1 U666 ( .A1(G111), .A2(n998), .ZN(n601) );
  NAND2_X1 U667 ( .A1(n602), .A2(n601), .ZN(n609) );
  NAND2_X1 U668 ( .A1(G123), .A2(n999), .ZN(n603) );
  XNOR2_X1 U669 ( .A(n603), .B(KEYINPUT18), .ZN(n607) );
  INV_X1 U670 ( .A(n604), .ZN(n605) );
  INV_X1 U671 ( .A(n605), .ZN(n1002) );
  NAND2_X1 U672 ( .A1(G135), .A2(n1002), .ZN(n606) );
  NAND2_X1 U673 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U674 ( .A1(n609), .A2(n608), .ZN(n986) );
  XNOR2_X1 U675 ( .A(n986), .B(G2096), .ZN(n611) );
  INV_X1 U676 ( .A(G2100), .ZN(n610) );
  NAND2_X1 U677 ( .A1(n611), .A2(n610), .ZN(G156) );
  NAND2_X1 U678 ( .A1(n907), .A2(G559), .ZN(n612) );
  XNOR2_X1 U679 ( .A(n612), .B(n1020), .ZN(n663) );
  NOR2_X1 U680 ( .A1(n663), .A2(G860), .ZN(n621) );
  NAND2_X1 U681 ( .A1(G80), .A2(n651), .ZN(n614) );
  NAND2_X1 U682 ( .A1(G93), .A2(n647), .ZN(n613) );
  NAND2_X1 U683 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U684 ( .A(KEYINPUT80), .B(n615), .ZN(n620) );
  NAND2_X1 U685 ( .A1(G55), .A2(n645), .ZN(n617) );
  NAND2_X1 U686 ( .A1(G67), .A2(n648), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n617), .A2(n616), .ZN(n618) );
  XOR2_X1 U688 ( .A(KEYINPUT81), .B(n618), .Z(n619) );
  OR2_X1 U689 ( .A1(n620), .A2(n619), .ZN(n667) );
  XOR2_X1 U690 ( .A(n621), .B(n667), .Z(G145) );
  NAND2_X1 U691 ( .A1(G49), .A2(n645), .ZN(n624) );
  NAND2_X1 U692 ( .A1(G87), .A2(n622), .ZN(n623) );
  NAND2_X1 U693 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U694 ( .A1(n648), .A2(n625), .ZN(n627) );
  NAND2_X1 U695 ( .A1(G651), .A2(G74), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n627), .A2(n626), .ZN(G288) );
  NAND2_X1 U697 ( .A1(n645), .A2(G47), .ZN(n634) );
  NAND2_X1 U698 ( .A1(G72), .A2(n651), .ZN(n629) );
  NAND2_X1 U699 ( .A1(G85), .A2(n647), .ZN(n628) );
  NAND2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U701 ( .A1(G60), .A2(n648), .ZN(n630) );
  XOR2_X1 U702 ( .A(KEYINPUT70), .B(n630), .Z(n631) );
  NOR2_X1 U703 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U704 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U705 ( .A(KEYINPUT71), .B(n635), .Z(G290) );
  NAND2_X1 U706 ( .A1(n647), .A2(G88), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n636), .B(KEYINPUT84), .ZN(n638) );
  NAND2_X1 U708 ( .A1(G75), .A2(n651), .ZN(n637) );
  NAND2_X1 U709 ( .A1(n638), .A2(n637), .ZN(n639) );
  XNOR2_X1 U710 ( .A(KEYINPUT85), .B(n639), .ZN(n644) );
  NAND2_X1 U711 ( .A1(G50), .A2(n645), .ZN(n641) );
  NAND2_X1 U712 ( .A1(G62), .A2(n648), .ZN(n640) );
  NAND2_X1 U713 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U714 ( .A(KEYINPUT83), .B(n642), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n644), .A2(n643), .ZN(G303) );
  INV_X1 U716 ( .A(G303), .ZN(G166) );
  NAND2_X1 U717 ( .A1(G48), .A2(n645), .ZN(n646) );
  XNOR2_X1 U718 ( .A(n646), .B(KEYINPUT82), .ZN(n656) );
  NAND2_X1 U719 ( .A1(G86), .A2(n647), .ZN(n650) );
  NAND2_X1 U720 ( .A1(G61), .A2(n648), .ZN(n649) );
  NAND2_X1 U721 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U722 ( .A1(n651), .A2(G73), .ZN(n652) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n652), .Z(n653) );
  NOR2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U725 ( .A1(n656), .A2(n655), .ZN(G305) );
  XOR2_X1 U726 ( .A(KEYINPUT86), .B(KEYINPUT19), .Z(n657) );
  XNOR2_X1 U727 ( .A(G288), .B(n657), .ZN(n658) );
  XOR2_X1 U728 ( .A(n667), .B(n658), .Z(n660) );
  XNOR2_X1 U729 ( .A(G290), .B(G166), .ZN(n659) );
  XNOR2_X1 U730 ( .A(n660), .B(n659), .ZN(n661) );
  INV_X1 U731 ( .A(G299), .ZN(n726) );
  XNOR2_X1 U732 ( .A(n661), .B(n726), .ZN(n662) );
  XNOR2_X1 U733 ( .A(n662), .B(G305), .ZN(n1016) );
  XNOR2_X1 U734 ( .A(n1016), .B(KEYINPUT87), .ZN(n664) );
  XNOR2_X1 U735 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U736 ( .A1(n665), .A2(G868), .ZN(n666) );
  XNOR2_X1 U737 ( .A(n666), .B(KEYINPUT88), .ZN(n670) );
  NAND2_X1 U738 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U739 ( .A1(n670), .A2(n669), .ZN(G295) );
  NAND2_X1 U740 ( .A1(G2078), .A2(G2084), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n671), .B(KEYINPUT20), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n672), .B(KEYINPUT89), .ZN(n673) );
  NAND2_X1 U743 ( .A1(n673), .A2(G2090), .ZN(n674) );
  XNOR2_X1 U744 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U745 ( .A1(n675), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U746 ( .A(KEYINPUT75), .B(G57), .ZN(G237) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U748 ( .A1(G237), .A2(G236), .ZN(n676) );
  NAND2_X1 U749 ( .A1(G69), .A2(n676), .ZN(n677) );
  XNOR2_X1 U750 ( .A(KEYINPUT91), .B(n677), .ZN(n678) );
  NAND2_X1 U751 ( .A1(n678), .A2(G108), .ZN(n964) );
  NAND2_X1 U752 ( .A1(n964), .A2(G567), .ZN(n684) );
  NAND2_X1 U753 ( .A1(G132), .A2(G82), .ZN(n679) );
  XNOR2_X1 U754 ( .A(n679), .B(KEYINPUT90), .ZN(n680) );
  XNOR2_X1 U755 ( .A(n680), .B(KEYINPUT22), .ZN(n681) );
  NOR2_X1 U756 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U757 ( .A1(G96), .A2(n682), .ZN(n965) );
  NAND2_X1 U758 ( .A1(n965), .A2(G2106), .ZN(n683) );
  NAND2_X1 U759 ( .A1(n684), .A2(n683), .ZN(n966) );
  NAND2_X1 U760 ( .A1(G483), .A2(G661), .ZN(n685) );
  NOR2_X1 U761 ( .A1(n966), .A2(n685), .ZN(n838) );
  NAND2_X1 U762 ( .A1(n838), .A2(G36), .ZN(n686) );
  XNOR2_X1 U763 ( .A(KEYINPUT92), .B(n686), .ZN(G176) );
  NAND2_X1 U764 ( .A1(G102), .A2(n1004), .ZN(n688) );
  NAND2_X1 U765 ( .A1(G138), .A2(n1002), .ZN(n687) );
  NAND2_X1 U766 ( .A1(n688), .A2(n687), .ZN(n692) );
  NAND2_X1 U767 ( .A1(G114), .A2(n998), .ZN(n690) );
  NAND2_X1 U768 ( .A1(G126), .A2(n999), .ZN(n689) );
  NAND2_X1 U769 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U770 ( .A1(n692), .A2(n691), .ZN(G164) );
  NAND2_X1 U771 ( .A1(G40), .A2(G160), .ZN(n781) );
  INV_X1 U772 ( .A(n781), .ZN(n693) );
  NOR2_X1 U773 ( .A1(G164), .A2(G1384), .ZN(n782) );
  NAND2_X2 U774 ( .A1(n693), .A2(n782), .ZN(n739) );
  NAND2_X1 U775 ( .A1(G8), .A2(n739), .ZN(n771) );
  NOR2_X1 U776 ( .A1(G1981), .A2(G305), .ZN(n694) );
  XOR2_X1 U777 ( .A(n694), .B(KEYINPUT24), .Z(n695) );
  NOR2_X1 U778 ( .A1(n771), .A2(n695), .ZN(n779) );
  NOR2_X1 U779 ( .A1(G2084), .A2(n739), .ZN(n696) );
  NAND2_X1 U780 ( .A1(G8), .A2(n696), .ZN(n738) );
  NOR2_X1 U781 ( .A1(G1966), .A2(n771), .ZN(n735) );
  NOR2_X1 U782 ( .A1(n735), .A2(n696), .ZN(n697) );
  NAND2_X1 U783 ( .A1(G8), .A2(n697), .ZN(n698) );
  XNOR2_X1 U784 ( .A(n698), .B(KEYINPUT30), .ZN(n699) );
  NOR2_X1 U785 ( .A1(n699), .A2(G168), .ZN(n703) );
  XNOR2_X1 U786 ( .A(G2078), .B(KEYINPUT25), .ZN(n888) );
  NOR2_X1 U787 ( .A1(n739), .A2(n888), .ZN(n701) );
  INV_X1 U788 ( .A(n739), .ZN(n708) );
  XNOR2_X1 U789 ( .A(G1961), .B(KEYINPUT97), .ZN(n931) );
  NOR2_X1 U790 ( .A1(n708), .A2(n931), .ZN(n700) );
  NOR2_X1 U791 ( .A1(n701), .A2(n700), .ZN(n706) );
  NOR2_X1 U792 ( .A1(G171), .A2(n706), .ZN(n702) );
  NOR2_X1 U793 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U794 ( .A(n704), .B(KEYINPUT31), .ZN(n705) );
  XNOR2_X1 U795 ( .A(n705), .B(KEYINPUT99), .ZN(n747) );
  NAND2_X1 U796 ( .A1(G171), .A2(n706), .ZN(n734) );
  NAND2_X1 U797 ( .A1(n708), .A2(G2072), .ZN(n707) );
  XNOR2_X1 U798 ( .A(n707), .B(KEYINPUT27), .ZN(n710) );
  INV_X1 U799 ( .A(G1956), .ZN(n942) );
  NOR2_X1 U800 ( .A1(n942), .A2(n708), .ZN(n709) );
  NOR2_X1 U801 ( .A1(n710), .A2(n709), .ZN(n727) );
  NOR2_X1 U802 ( .A1(n727), .A2(n726), .ZN(n712) );
  INV_X1 U803 ( .A(KEYINPUT28), .ZN(n711) );
  XNOR2_X1 U804 ( .A(n712), .B(n711), .ZN(n731) );
  INV_X1 U805 ( .A(G1996), .ZN(n889) );
  INV_X1 U806 ( .A(KEYINPUT26), .ZN(n713) );
  XNOR2_X1 U807 ( .A(n714), .B(n713), .ZN(n717) );
  AND2_X1 U808 ( .A1(n739), .A2(G1341), .ZN(n715) );
  NOR2_X1 U809 ( .A1(n715), .A2(n1020), .ZN(n716) );
  AND2_X1 U810 ( .A1(n717), .A2(n716), .ZN(n723) );
  NAND2_X1 U811 ( .A1(n723), .A2(n907), .ZN(n722) );
  INV_X1 U812 ( .A(G2067), .ZN(n886) );
  NOR2_X1 U813 ( .A1(n739), .A2(n886), .ZN(n718) );
  XOR2_X1 U814 ( .A(n718), .B(KEYINPUT98), .Z(n720) );
  NAND2_X1 U815 ( .A1(n739), .A2(G1348), .ZN(n719) );
  NAND2_X1 U816 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U817 ( .A1(n722), .A2(n721), .ZN(n725) );
  OR2_X1 U818 ( .A1(n907), .A2(n723), .ZN(n724) );
  NAND2_X1 U819 ( .A1(n725), .A2(n724), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n727), .A2(n726), .ZN(n728) );
  NAND2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U822 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U823 ( .A(n732), .B(KEYINPUT29), .Z(n733) );
  NAND2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n745) );
  AND2_X1 U825 ( .A1(n747), .A2(n745), .ZN(n736) );
  NOR2_X1 U826 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U827 ( .A1(n738), .A2(n737), .ZN(n754) );
  INV_X1 U828 ( .A(G8), .ZN(n744) );
  NOR2_X1 U829 ( .A1(G1971), .A2(n771), .ZN(n741) );
  NOR2_X1 U830 ( .A1(G2090), .A2(n739), .ZN(n740) );
  NOR2_X1 U831 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U832 ( .A1(n742), .A2(G303), .ZN(n743) );
  OR2_X1 U833 ( .A1(n744), .A2(n743), .ZN(n748) );
  AND2_X1 U834 ( .A1(n745), .A2(n748), .ZN(n746) );
  NAND2_X1 U835 ( .A1(n747), .A2(n746), .ZN(n751) );
  INV_X1 U836 ( .A(n748), .ZN(n749) );
  OR2_X1 U837 ( .A1(n749), .A2(G286), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U839 ( .A(n752), .B(KEYINPUT32), .ZN(n753) );
  NAND2_X1 U840 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U841 ( .A(KEYINPUT100), .B(n755), .ZN(n764) );
  NAND2_X1 U842 ( .A1(G166), .A2(G8), .ZN(n756) );
  OR2_X1 U843 ( .A1(G2090), .A2(n756), .ZN(n757) );
  AND2_X1 U844 ( .A1(n764), .A2(n757), .ZN(n759) );
  INV_X1 U845 ( .A(KEYINPUT102), .ZN(n758) );
  XNOR2_X1 U846 ( .A(n759), .B(n758), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n760), .A2(n771), .ZN(n777) );
  NOR2_X1 U848 ( .A1(G1976), .A2(G288), .ZN(n770) );
  NOR2_X1 U849 ( .A1(G1971), .A2(G303), .ZN(n761) );
  NOR2_X1 U850 ( .A1(n770), .A2(n761), .ZN(n915) );
  INV_X1 U851 ( .A(KEYINPUT33), .ZN(n762) );
  AND2_X1 U852 ( .A1(n915), .A2(n762), .ZN(n763) );
  NAND2_X1 U853 ( .A1(n764), .A2(n763), .ZN(n769) );
  NAND2_X1 U854 ( .A1(G288), .A2(G1976), .ZN(n765) );
  XOR2_X1 U855 ( .A(KEYINPUT101), .B(n765), .Z(n911) );
  INV_X1 U856 ( .A(n911), .ZN(n766) );
  NOR2_X1 U857 ( .A1(n766), .A2(n771), .ZN(n767) );
  OR2_X1 U858 ( .A1(KEYINPUT33), .A2(n767), .ZN(n768) );
  NAND2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n774) );
  NAND2_X1 U860 ( .A1(n770), .A2(KEYINPUT33), .ZN(n772) );
  NOR2_X1 U861 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U862 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U863 ( .A(G1981), .B(G305), .Z(n921) );
  NAND2_X1 U864 ( .A1(n775), .A2(n921), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U866 ( .A(n780), .B(KEYINPUT103), .ZN(n816) );
  XNOR2_X1 U867 ( .A(G1986), .B(G290), .ZN(n917) );
  NOR2_X1 U868 ( .A1(n782), .A2(n781), .ZN(n829) );
  NAND2_X1 U869 ( .A1(n917), .A2(n829), .ZN(n814) );
  INV_X1 U870 ( .A(G1991), .ZN(n818) );
  NAND2_X1 U871 ( .A1(G119), .A2(n999), .ZN(n789) );
  NAND2_X1 U872 ( .A1(G95), .A2(n1004), .ZN(n784) );
  NAND2_X1 U873 ( .A1(G107), .A2(n998), .ZN(n783) );
  NAND2_X1 U874 ( .A1(n784), .A2(n783), .ZN(n787) );
  NAND2_X1 U875 ( .A1(G131), .A2(n1002), .ZN(n785) );
  XNOR2_X1 U876 ( .A(KEYINPUT95), .B(n785), .ZN(n786) );
  NOR2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U879 ( .A(n790), .B(KEYINPUT96), .Z(n994) );
  NOR2_X1 U880 ( .A1(n818), .A2(n994), .ZN(n799) );
  NAND2_X1 U881 ( .A1(G117), .A2(n998), .ZN(n792) );
  NAND2_X1 U882 ( .A1(G129), .A2(n999), .ZN(n791) );
  NAND2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n1004), .A2(G105), .ZN(n793) );
  XOR2_X1 U885 ( .A(KEYINPUT38), .B(n793), .Z(n794) );
  NOR2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n797) );
  NAND2_X1 U887 ( .A1(G141), .A2(n1002), .ZN(n796) );
  NAND2_X1 U888 ( .A1(n797), .A2(n796), .ZN(n988) );
  AND2_X1 U889 ( .A1(G1996), .A2(n988), .ZN(n798) );
  NOR2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n848) );
  INV_X1 U891 ( .A(n829), .ZN(n800) );
  NOR2_X1 U892 ( .A1(n848), .A2(n800), .ZN(n821) );
  NAND2_X1 U893 ( .A1(G104), .A2(n1004), .ZN(n802) );
  NAND2_X1 U894 ( .A1(G140), .A2(n1002), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U896 ( .A(KEYINPUT34), .B(n803), .ZN(n809) );
  NAND2_X1 U897 ( .A1(G116), .A2(n998), .ZN(n805) );
  NAND2_X1 U898 ( .A1(G128), .A2(n999), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n806) );
  XNOR2_X1 U900 ( .A(KEYINPUT35), .B(n806), .ZN(n807) );
  XNOR2_X1 U901 ( .A(KEYINPUT93), .B(n807), .ZN(n808) );
  NOR2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n810) );
  XNOR2_X1 U903 ( .A(KEYINPUT36), .B(n810), .ZN(n995) );
  XNOR2_X1 U904 ( .A(G2067), .B(KEYINPUT37), .ZN(n826) );
  NOR2_X1 U905 ( .A1(n995), .A2(n826), .ZN(n876) );
  NAND2_X1 U906 ( .A1(n876), .A2(n829), .ZN(n811) );
  XNOR2_X1 U907 ( .A(n811), .B(KEYINPUT94), .ZN(n824) );
  INV_X1 U908 ( .A(n824), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n821), .A2(n812), .ZN(n813) );
  AND2_X1 U910 ( .A1(n814), .A2(n813), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n816), .A2(n815), .ZN(n832) );
  NOR2_X1 U912 ( .A1(n988), .A2(G1996), .ZN(n817) );
  XNOR2_X1 U913 ( .A(n817), .B(KEYINPUT104), .ZN(n866) );
  NOR2_X1 U914 ( .A1(G1986), .A2(G290), .ZN(n819) );
  AND2_X1 U915 ( .A1(n818), .A2(n994), .ZN(n870) );
  NOR2_X1 U916 ( .A1(n819), .A2(n870), .ZN(n820) );
  NOR2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n822) );
  NOR2_X1 U918 ( .A1(n866), .A2(n822), .ZN(n823) );
  XNOR2_X1 U919 ( .A(KEYINPUT39), .B(n823), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n825), .A2(n824), .ZN(n827) );
  NAND2_X1 U921 ( .A1(n995), .A2(n826), .ZN(n847) );
  NAND2_X1 U922 ( .A1(n827), .A2(n847), .ZN(n828) );
  XOR2_X1 U923 ( .A(KEYINPUT105), .B(n828), .Z(n830) );
  NAND2_X1 U924 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n832), .A2(n831), .ZN(n834) );
  XNOR2_X1 U926 ( .A(KEYINPUT40), .B(KEYINPUT106), .ZN(n833) );
  XNOR2_X1 U927 ( .A(n834), .B(n833), .ZN(G329) );
  NAND2_X1 U928 ( .A1(G2106), .A2(n835), .ZN(G217) );
  AND2_X1 U929 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U930 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U931 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U932 ( .A1(n838), .A2(n837), .ZN(G188) );
  NAND2_X1 U934 ( .A1(G100), .A2(n1004), .ZN(n840) );
  NAND2_X1 U935 ( .A1(G112), .A2(n998), .ZN(n839) );
  NAND2_X1 U936 ( .A1(n840), .A2(n839), .ZN(n846) );
  NAND2_X1 U937 ( .A1(G124), .A2(n999), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n841), .B(KEYINPUT44), .ZN(n844) );
  NAND2_X1 U939 ( .A1(n1002), .A2(G136), .ZN(n842) );
  XNOR2_X1 U940 ( .A(n842), .B(KEYINPUT110), .ZN(n843) );
  NAND2_X1 U941 ( .A1(n844), .A2(n843), .ZN(n845) );
  NOR2_X1 U942 ( .A1(n846), .A2(n845), .ZN(G162) );
  NAND2_X1 U943 ( .A1(n848), .A2(n847), .ZN(n863) );
  NAND2_X1 U944 ( .A1(G103), .A2(n1004), .ZN(n850) );
  NAND2_X1 U945 ( .A1(G139), .A2(n1002), .ZN(n849) );
  NAND2_X1 U946 ( .A1(n850), .A2(n849), .ZN(n856) );
  NAND2_X1 U947 ( .A1(G115), .A2(n998), .ZN(n852) );
  NAND2_X1 U948 ( .A1(G127), .A2(n999), .ZN(n851) );
  NAND2_X1 U949 ( .A1(n852), .A2(n851), .ZN(n853) );
  XOR2_X1 U950 ( .A(KEYINPUT112), .B(n853), .Z(n854) );
  XNOR2_X1 U951 ( .A(KEYINPUT47), .B(n854), .ZN(n855) );
  NOR2_X1 U952 ( .A1(n856), .A2(n855), .ZN(n857) );
  XOR2_X1 U953 ( .A(KEYINPUT113), .B(n857), .Z(n987) );
  XOR2_X1 U954 ( .A(G2072), .B(n987), .Z(n859) );
  XOR2_X1 U955 ( .A(G164), .B(G2078), .Z(n858) );
  NOR2_X1 U956 ( .A1(n859), .A2(n858), .ZN(n860) );
  XOR2_X1 U957 ( .A(KEYINPUT50), .B(n860), .Z(n861) );
  XNOR2_X1 U958 ( .A(KEYINPUT120), .B(n861), .ZN(n862) );
  NOR2_X1 U959 ( .A1(n863), .A2(n862), .ZN(n869) );
  XNOR2_X1 U960 ( .A(G2090), .B(G162), .ZN(n864) );
  XNOR2_X1 U961 ( .A(n864), .B(KEYINPUT119), .ZN(n865) );
  NOR2_X1 U962 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U963 ( .A(KEYINPUT51), .B(n867), .Z(n868) );
  NAND2_X1 U964 ( .A1(n869), .A2(n868), .ZN(n879) );
  NOR2_X1 U965 ( .A1(n870), .A2(n986), .ZN(n871) );
  XOR2_X1 U966 ( .A(KEYINPUT116), .B(n871), .Z(n873) );
  XOR2_X1 U967 ( .A(G160), .B(G2084), .Z(n872) );
  NOR2_X1 U968 ( .A1(n873), .A2(n872), .ZN(n874) );
  XNOR2_X1 U969 ( .A(n874), .B(KEYINPUT117), .ZN(n875) );
  NOR2_X1 U970 ( .A1(n876), .A2(n875), .ZN(n877) );
  XOR2_X1 U971 ( .A(KEYINPUT118), .B(n877), .Z(n878) );
  NOR2_X1 U972 ( .A1(n879), .A2(n878), .ZN(n880) );
  XNOR2_X1 U973 ( .A(KEYINPUT52), .B(n880), .ZN(n882) );
  INV_X1 U974 ( .A(KEYINPUT55), .ZN(n881) );
  NAND2_X1 U975 ( .A1(n882), .A2(n881), .ZN(n883) );
  NAND2_X1 U976 ( .A1(n883), .A2(G29), .ZN(n962) );
  XNOR2_X1 U977 ( .A(G29), .B(KEYINPUT121), .ZN(n904) );
  XNOR2_X1 U978 ( .A(G1991), .B(G25), .ZN(n885) );
  XNOR2_X1 U979 ( .A(G33), .B(G2072), .ZN(n884) );
  NOR2_X1 U980 ( .A1(n885), .A2(n884), .ZN(n895) );
  XNOR2_X1 U981 ( .A(G26), .B(n886), .ZN(n887) );
  NAND2_X1 U982 ( .A1(n887), .A2(G28), .ZN(n893) );
  XNOR2_X1 U983 ( .A(n888), .B(G27), .ZN(n891) );
  XNOR2_X1 U984 ( .A(n889), .B(G32), .ZN(n890) );
  NAND2_X1 U985 ( .A1(n891), .A2(n890), .ZN(n892) );
  NOR2_X1 U986 ( .A1(n893), .A2(n892), .ZN(n894) );
  NAND2_X1 U987 ( .A1(n895), .A2(n894), .ZN(n896) );
  XNOR2_X1 U988 ( .A(n896), .B(KEYINPUT53), .ZN(n899) );
  XOR2_X1 U989 ( .A(G2084), .B(G34), .Z(n897) );
  XNOR2_X1 U990 ( .A(KEYINPUT54), .B(n897), .ZN(n898) );
  NAND2_X1 U991 ( .A1(n899), .A2(n898), .ZN(n901) );
  XNOR2_X1 U992 ( .A(G35), .B(G2090), .ZN(n900) );
  NOR2_X1 U993 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U994 ( .A(KEYINPUT55), .B(n902), .ZN(n903) );
  NAND2_X1 U995 ( .A1(n904), .A2(n903), .ZN(n905) );
  XNOR2_X1 U996 ( .A(KEYINPUT122), .B(n905), .ZN(n906) );
  NAND2_X1 U997 ( .A1(n906), .A2(G11), .ZN(n960) );
  XNOR2_X1 U998 ( .A(G16), .B(KEYINPUT56), .ZN(n930) );
  XNOR2_X1 U999 ( .A(G171), .B(G1961), .ZN(n909) );
  XNOR2_X1 U1000 ( .A(n907), .B(G1348), .ZN(n908) );
  NAND2_X1 U1001 ( .A1(n909), .A2(n908), .ZN(n920) );
  NAND2_X1 U1002 ( .A1(G1971), .A2(G303), .ZN(n910) );
  NAND2_X1 U1003 ( .A1(n911), .A2(n910), .ZN(n913) );
  XNOR2_X1 U1004 ( .A(G1956), .B(G299), .ZN(n912) );
  NOR2_X1 U1005 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1006 ( .A1(n915), .A2(n914), .ZN(n916) );
  NOR2_X1 U1007 ( .A1(n917), .A2(n916), .ZN(n918) );
  XOR2_X1 U1008 ( .A(KEYINPUT124), .B(n918), .Z(n919) );
  NOR2_X1 U1009 ( .A1(n920), .A2(n919), .ZN(n928) );
  XNOR2_X1 U1010 ( .A(n1020), .B(G1341), .ZN(n926) );
  XNOR2_X1 U1011 ( .A(G1966), .B(G168), .ZN(n922) );
  NAND2_X1 U1012 ( .A1(n922), .A2(n921), .ZN(n923) );
  XNOR2_X1 U1013 ( .A(n923), .B(KEYINPUT57), .ZN(n924) );
  XNOR2_X1 U1014 ( .A(KEYINPUT123), .B(n924), .ZN(n925) );
  NOR2_X1 U1015 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1016 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1017 ( .A1(n930), .A2(n929), .ZN(n958) );
  INV_X1 U1018 ( .A(G16), .ZN(n956) );
  XNOR2_X1 U1019 ( .A(KEYINPUT125), .B(G5), .ZN(n932) );
  XNOR2_X1 U1020 ( .A(n932), .B(n931), .ZN(n939) );
  XNOR2_X1 U1021 ( .A(G1971), .B(G22), .ZN(n934) );
  XNOR2_X1 U1022 ( .A(G23), .B(G1976), .ZN(n933) );
  NOR2_X1 U1023 ( .A1(n934), .A2(n933), .ZN(n936) );
  XOR2_X1 U1024 ( .A(G1986), .B(G24), .Z(n935) );
  NAND2_X1 U1025 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1026 ( .A(KEYINPUT58), .B(n937), .ZN(n938) );
  NOR2_X1 U1027 ( .A1(n939), .A2(n938), .ZN(n951) );
  XOR2_X1 U1028 ( .A(G4), .B(KEYINPUT126), .Z(n941) );
  XNOR2_X1 U1029 ( .A(G1348), .B(KEYINPUT59), .ZN(n940) );
  XNOR2_X1 U1030 ( .A(n941), .B(n940), .ZN(n948) );
  XNOR2_X1 U1031 ( .A(G20), .B(n942), .ZN(n946) );
  XNOR2_X1 U1032 ( .A(G1341), .B(G19), .ZN(n944) );
  XNOR2_X1 U1033 ( .A(G1981), .B(G6), .ZN(n943) );
  NOR2_X1 U1034 ( .A1(n944), .A2(n943), .ZN(n945) );
  NAND2_X1 U1035 ( .A1(n946), .A2(n945), .ZN(n947) );
  NOR2_X1 U1036 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1037 ( .A(n949), .B(KEYINPUT60), .ZN(n950) );
  NAND2_X1 U1038 ( .A1(n951), .A2(n950), .ZN(n953) );
  XNOR2_X1 U1039 ( .A(G21), .B(G1966), .ZN(n952) );
  NOR2_X1 U1040 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1041 ( .A(KEYINPUT61), .B(n954), .ZN(n955) );
  NAND2_X1 U1042 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1043 ( .A1(n958), .A2(n957), .ZN(n959) );
  NOR2_X1 U1044 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1045 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1046 ( .A(KEYINPUT62), .B(n963), .Z(G311) );
  XNOR2_X1 U1047 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
  INV_X1 U1048 ( .A(G132), .ZN(G219) );
  INV_X1 U1049 ( .A(G108), .ZN(G238) );
  INV_X1 U1050 ( .A(G82), .ZN(G220) );
  NOR2_X1 U1051 ( .A1(n965), .A2(n964), .ZN(G325) );
  INV_X1 U1052 ( .A(G325), .ZN(G261) );
  INV_X1 U1053 ( .A(n966), .ZN(G319) );
  XOR2_X1 U1054 ( .A(KEYINPUT109), .B(G2678), .Z(n968) );
  XNOR2_X1 U1055 ( .A(G2072), .B(G2090), .ZN(n967) );
  XNOR2_X1 U1056 ( .A(n968), .B(n967), .ZN(n972) );
  XOR2_X1 U1057 ( .A(KEYINPUT43), .B(KEYINPUT108), .Z(n970) );
  XNOR2_X1 U1058 ( .A(G2067), .B(KEYINPUT42), .ZN(n969) );
  XNOR2_X1 U1059 ( .A(n970), .B(n969), .ZN(n971) );
  XOR2_X1 U1060 ( .A(n972), .B(n971), .Z(n974) );
  XNOR2_X1 U1061 ( .A(G2096), .B(G2100), .ZN(n973) );
  XNOR2_X1 U1062 ( .A(n974), .B(n973), .ZN(n976) );
  XOR2_X1 U1063 ( .A(G2078), .B(G2084), .Z(n975) );
  XNOR2_X1 U1064 ( .A(n976), .B(n975), .ZN(G227) );
  XOR2_X1 U1065 ( .A(G1976), .B(G1981), .Z(n978) );
  XNOR2_X1 U1066 ( .A(G1966), .B(G1971), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(n978), .B(n977), .ZN(n979) );
  XOR2_X1 U1068 ( .A(n979), .B(KEYINPUT41), .Z(n981) );
  XNOR2_X1 U1069 ( .A(G1991), .B(G2474), .ZN(n980) );
  XNOR2_X1 U1070 ( .A(n981), .B(n980), .ZN(n985) );
  XOR2_X1 U1071 ( .A(G1956), .B(G1961), .Z(n983) );
  XNOR2_X1 U1072 ( .A(G1996), .B(G1986), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(n983), .B(n982), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(n985), .B(n984), .ZN(G229) );
  XNOR2_X1 U1075 ( .A(n987), .B(n986), .ZN(n990) );
  XOR2_X1 U1076 ( .A(G160), .B(n988), .Z(n989) );
  XNOR2_X1 U1077 ( .A(n990), .B(n989), .ZN(n1013) );
  XOR2_X1 U1078 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n992) );
  XNOR2_X1 U1079 ( .A(G164), .B(KEYINPUT46), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(n992), .B(n991), .ZN(n993) );
  XNOR2_X1 U1081 ( .A(G162), .B(n993), .ZN(n997) );
  XOR2_X1 U1082 ( .A(n995), .B(n994), .Z(n996) );
  XNOR2_X1 U1083 ( .A(n997), .B(n996), .ZN(n1011) );
  NAND2_X1 U1084 ( .A1(G118), .A2(n998), .ZN(n1001) );
  NAND2_X1 U1085 ( .A1(G130), .A2(n999), .ZN(n1000) );
  NAND2_X1 U1086 ( .A1(n1001), .A2(n1000), .ZN(n1009) );
  NAND2_X1 U1087 ( .A1(G142), .A2(n1002), .ZN(n1003) );
  XOR2_X1 U1088 ( .A(KEYINPUT111), .B(n1003), .Z(n1006) );
  NAND2_X1 U1089 ( .A1(n1004), .A2(G106), .ZN(n1005) );
  NAND2_X1 U1090 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1091 ( .A(n1007), .B(KEYINPUT45), .Z(n1008) );
  NOR2_X1 U1092 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1093 ( .A(n1011), .B(n1010), .Z(n1012) );
  XOR2_X1 U1094 ( .A(n1013), .B(n1012), .Z(n1014) );
  NOR2_X1 U1095 ( .A1(G37), .A2(n1014), .ZN(n1015) );
  XOR2_X1 U1096 ( .A(KEYINPUT115), .B(n1015), .Z(G395) );
  XOR2_X1 U1097 ( .A(n1016), .B(G286), .Z(n1019) );
  XNOR2_X1 U1098 ( .A(G171), .B(n1017), .ZN(n1018) );
  XNOR2_X1 U1099 ( .A(n1019), .B(n1018), .ZN(n1021) );
  XNOR2_X1 U1100 ( .A(n1021), .B(n1020), .ZN(n1022) );
  NOR2_X1 U1101 ( .A1(G37), .A2(n1022), .ZN(G397) );
  XOR2_X1 U1102 ( .A(G2443), .B(G2454), .Z(n1024) );
  XNOR2_X1 U1103 ( .A(G1348), .B(G2435), .ZN(n1023) );
  XNOR2_X1 U1104 ( .A(n1024), .B(n1023), .ZN(n1031) );
  XOR2_X1 U1105 ( .A(KEYINPUT107), .B(G2446), .Z(n1026) );
  XNOR2_X1 U1106 ( .A(G1341), .B(G2430), .ZN(n1025) );
  XNOR2_X1 U1107 ( .A(n1026), .B(n1025), .ZN(n1027) );
  XOR2_X1 U1108 ( .A(n1027), .B(G2451), .Z(n1029) );
  XNOR2_X1 U1109 ( .A(G2438), .B(G2427), .ZN(n1028) );
  XNOR2_X1 U1110 ( .A(n1029), .B(n1028), .ZN(n1030) );
  XNOR2_X1 U1111 ( .A(n1031), .B(n1030), .ZN(n1032) );
  NAND2_X1 U1112 ( .A1(n1032), .A2(G14), .ZN(n1038) );
  NAND2_X1 U1113 ( .A1(G319), .A2(n1038), .ZN(n1035) );
  NOR2_X1 U1114 ( .A1(G227), .A2(G229), .ZN(n1033) );
  XNOR2_X1 U1115 ( .A(KEYINPUT49), .B(n1033), .ZN(n1034) );
  NOR2_X1 U1116 ( .A1(n1035), .A2(n1034), .ZN(n1037) );
  NOR2_X1 U1117 ( .A1(G395), .A2(G397), .ZN(n1036) );
  NAND2_X1 U1118 ( .A1(n1037), .A2(n1036), .ZN(G225) );
  INV_X1 U1119 ( .A(G225), .ZN(G308) );
  INV_X1 U1120 ( .A(G96), .ZN(G221) );
  INV_X1 U1121 ( .A(G69), .ZN(G235) );
  INV_X1 U1122 ( .A(n1038), .ZN(G401) );
endmodule

