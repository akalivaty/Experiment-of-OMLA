//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:00 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G140), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G125), .ZN(new_n193));
  INV_X1    g007(.A(G125), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G140), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT74), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n192), .A2(KEYINPUT74), .A3(G125), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(KEYINPUT16), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT16), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n193), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n199), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n199), .A2(new_n204), .A3(new_n201), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G110), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT73), .ZN(new_n208));
  XNOR2_X1  g022(.A(KEYINPUT67), .B(G119), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G128), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT67), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT67), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G119), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n212), .A2(new_n214), .A3(G128), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(KEYINPUT23), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n212), .A2(new_n214), .ZN(new_n217));
  INV_X1    g031(.A(G128), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(KEYINPUT73), .A3(new_n218), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n210), .A2(new_n216), .A3(new_n219), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(KEYINPUT23), .A3(G119), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n207), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n215), .B1(new_n211), .B2(G128), .ZN(new_n223));
  XNOR2_X1  g037(.A(KEYINPUT24), .B(G110), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n206), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  AND2_X1   g040(.A1(new_n193), .A2(new_n195), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n204), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n203), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n220), .A2(new_n207), .A3(new_n221), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n223), .A2(new_n224), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n191), .B1(new_n226), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n222), .A2(new_n225), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n203), .A2(new_n205), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n230), .A2(new_n231), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(new_n203), .A3(new_n228), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n238), .A3(new_n190), .ZN(new_n239));
  INV_X1    g053(.A(G217), .ZN(new_n240));
  INV_X1    g054(.A(G902), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n240), .B1(G234), .B2(new_n241), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n242), .A2(G902), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n233), .A2(new_n239), .A3(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n233), .A2(new_n241), .A3(new_n239), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT25), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n233), .A2(KEYINPUT25), .A3(new_n239), .A4(new_n241), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n244), .B1(new_n249), .B2(new_n242), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(G472), .A2(G902), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT70), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT68), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n204), .A2(G143), .ZN(new_n256));
  INV_X1    g070(.A(G143), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G146), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n255), .A2(new_n256), .A3(new_n258), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT1), .B1(new_n257), .B2(G146), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT66), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g076(.A(KEYINPUT66), .B(KEYINPUT1), .C1(new_n257), .C2(G146), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(G128), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n256), .A2(new_n258), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n259), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G137), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT65), .A3(G134), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n269));
  INV_X1    g083(.A(G134), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n269), .B1(new_n270), .B2(G137), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n267), .A2(G134), .ZN(new_n272));
  OAI211_X1 g086(.A(G131), .B(new_n268), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT11), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n274), .B1(new_n270), .B2(G137), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n267), .A2(KEYINPUT11), .A3(G134), .ZN(new_n276));
  INV_X1    g090(.A(G131), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n270), .A2(G137), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n275), .A2(new_n276), .A3(new_n277), .A4(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n254), .B1(new_n266), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n263), .A2(G128), .ZN(new_n282));
  AOI21_X1  g096(.A(KEYINPUT66), .B1(new_n256), .B2(KEYINPUT1), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n265), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n259), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n280), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(KEYINPUT68), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n275), .A2(new_n276), .A3(new_n278), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G131), .ZN(new_n290));
  OR2_X1    g104(.A1(KEYINPUT0), .A2(G128), .ZN(new_n291));
  NAND2_X1  g105(.A1(KEYINPUT0), .A2(G128), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n265), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n256), .A2(new_n258), .A3(new_n292), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n290), .A2(new_n279), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n281), .A2(new_n288), .A3(KEYINPUT30), .A4(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT30), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n290), .A2(new_n279), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT64), .ZN(new_n301));
  AOI22_X1  g115(.A1(new_n256), .A2(new_n258), .B1(new_n291), .B2(new_n292), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n256), .A2(new_n258), .A3(new_n292), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n294), .A2(KEYINPUT64), .A3(new_n295), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n300), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n280), .B1(new_n285), .B2(new_n284), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n299), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n212), .A2(new_n214), .A3(G116), .ZN(new_n309));
  INV_X1    g123(.A(G116), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G119), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT2), .B(G113), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n313), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n315), .A2(new_n309), .A3(new_n311), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n298), .A2(new_n308), .A3(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(new_n314), .A2(new_n316), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n281), .A2(new_n288), .A3(new_n297), .A4(new_n319), .ZN(new_n320));
  XOR2_X1   g134(.A(KEYINPUT26), .B(G101), .Z(new_n321));
  NOR2_X1   g135(.A1(G237), .A2(G953), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G210), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n321), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n320), .A2(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(new_n253), .B1(new_n318), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n286), .A2(new_n287), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n300), .A2(new_n304), .A3(new_n305), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n319), .B1(new_n331), .B2(new_n299), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n298), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n333), .A2(KEYINPUT70), .A3(new_n320), .A4(new_n326), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n328), .A2(KEYINPUT31), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n327), .B1(new_n298), .B2(new_n332), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT31), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT28), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n331), .A2(new_n317), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(new_n320), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n329), .A2(new_n297), .A3(new_n319), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT71), .B1(new_n342), .B2(new_n339), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT71), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n317), .A2(new_n296), .ZN(new_n345));
  AOI211_X1 g159(.A(new_n344), .B(KEYINPUT28), .C1(new_n345), .C2(new_n329), .ZN(new_n346));
  NOR3_X1   g160(.A1(new_n341), .A2(new_n343), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n338), .B1(new_n326), .B2(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n252), .B1(new_n335), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT32), .ZN(new_n350));
  INV_X1    g164(.A(new_n252), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n346), .A2(new_n343), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n340), .A2(new_n320), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT28), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(new_n326), .ZN(new_n356));
  AOI22_X1  g170(.A1(new_n355), .A2(new_n356), .B1(new_n336), .B2(new_n337), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n328), .A2(KEYINPUT31), .A3(new_n334), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n351), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT32), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n350), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT72), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n346), .B2(new_n343), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n296), .B1(new_n307), .B2(KEYINPUT68), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n319), .B1(new_n365), .B2(new_n281), .ZN(new_n366));
  AND4_X1   g180(.A1(new_n281), .A2(new_n288), .A3(new_n297), .A4(new_n319), .ZN(new_n367));
  OAI21_X1  g181(.A(KEYINPUT28), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n307), .A2(new_n296), .A3(new_n317), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n344), .B1(new_n369), .B2(KEYINPUT28), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n342), .A2(KEYINPUT71), .A3(new_n339), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(KEYINPUT72), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT29), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n356), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n364), .A2(new_n368), .A3(new_n372), .A4(new_n374), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n375), .A2(new_n241), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n333), .A2(new_n320), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n356), .ZN(new_n378));
  OAI211_X1 g192(.A(new_n378), .B(new_n373), .C1(new_n355), .C2(new_n356), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G472), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n251), .B1(new_n362), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G469), .ZN(new_n383));
  XNOR2_X1  g197(.A(G110), .B(G140), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n188), .A2(G227), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n384), .B(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G104), .ZN(new_n387));
  OAI21_X1  g201(.A(KEYINPUT3), .B1(new_n387), .B2(G107), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(G104), .ZN(new_n391));
  INV_X1    g205(.A(G101), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n387), .A2(G107), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n388), .A2(new_n391), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n387), .A2(G107), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n390), .A2(G104), .ZN(new_n396));
  OAI21_X1  g210(.A(G101), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n394), .A2(new_n397), .A3(KEYINPUT10), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n286), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n294), .A2(new_n295), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n388), .A2(new_n391), .A3(new_n393), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n401), .A2(new_n402), .A3(G101), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n401), .A2(G101), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n394), .A2(KEYINPUT4), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n400), .B(new_n403), .C1(new_n404), .C2(new_n405), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n260), .A2(G128), .B1(new_n256), .B2(new_n258), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n397), .B(new_n394), .C1(new_n407), .C2(new_n259), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT10), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n399), .A2(new_n406), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT77), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n399), .A2(new_n406), .A3(new_n410), .A4(KEYINPUT77), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n413), .A2(new_n300), .A3(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n300), .B(KEYINPUT75), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n386), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n386), .B1(new_n411), .B2(new_n416), .ZN(new_n420));
  INV_X1    g234(.A(new_n300), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n394), .A2(new_n397), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n284), .A2(new_n422), .A3(new_n285), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n421), .B1(new_n423), .B2(new_n408), .ZN(new_n424));
  AOI21_X1  g238(.A(KEYINPUT12), .B1(new_n300), .B2(KEYINPUT76), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(new_n426), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n420), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n383), .B(new_n241), .C1(new_n419), .C2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT78), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n421), .B1(new_n411), .B2(new_n412), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n417), .B1(new_n433), .B2(new_n414), .ZN(new_n434));
  INV_X1    g248(.A(new_n429), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(new_n427), .ZN(new_n436));
  OAI22_X1  g250(.A1(new_n434), .A2(new_n386), .B1(new_n436), .B2(new_n420), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT78), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n437), .A2(new_n438), .A3(new_n383), .A4(new_n241), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n432), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n420), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n415), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n417), .B1(new_n429), .B2(new_n428), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(new_n386), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n383), .B1(new_n444), .B2(new_n241), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G210), .B1(G237), .B2(G902), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(KEYINPUT81), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT80), .B(G224), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(G953), .ZN(new_n451));
  AOI21_X1  g265(.A(G125), .B1(new_n284), .B2(new_n285), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n194), .B1(new_n294), .B2(new_n295), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n453), .ZN(new_n455));
  INV_X1    g269(.A(new_n451), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n455), .B(new_n456), .C1(new_n266), .C2(G125), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n401), .A2(G101), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n459), .A2(KEYINPUT4), .A3(new_n394), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n317), .A2(new_n460), .A3(new_n403), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT5), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n209), .A2(new_n462), .A3(G116), .ZN(new_n463));
  OAI211_X1 g277(.A(G113), .B(new_n463), .C1(new_n312), .C2(new_n462), .ZN(new_n464));
  INV_X1    g278(.A(new_n422), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n464), .A2(new_n316), .A3(new_n465), .ZN(new_n466));
  XNOR2_X1  g280(.A(G110), .B(G122), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n461), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT6), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n461), .A2(new_n466), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT79), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(KEYINPUT6), .A3(new_n472), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n458), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT7), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n456), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n454), .A2(new_n457), .A3(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(new_n467), .B(KEYINPUT8), .ZN(new_n480));
  AND3_X1   g294(.A1(new_n464), .A2(new_n316), .A3(new_n465), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n465), .B1(new_n464), .B2(new_n316), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n452), .A2(new_n453), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n484), .A2(new_n477), .A3(new_n456), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n479), .A2(new_n483), .A3(new_n468), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n241), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n449), .B1(new_n476), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(new_n458), .ZN(new_n489));
  AOI22_X1  g303(.A1(new_n468), .A2(KEYINPUT6), .B1(new_n470), .B2(new_n472), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n470), .A2(KEYINPUT6), .A3(new_n472), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(new_n241), .A3(new_n448), .A4(new_n486), .ZN(new_n493));
  AND2_X1   g307(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G214), .B1(G237), .B2(G902), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT9), .B(G234), .ZN(new_n498));
  OAI21_X1  g312(.A(G221), .B1(new_n498), .B2(G902), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n447), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT85), .ZN(new_n501));
  XNOR2_X1  g315(.A(G113), .B(G122), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(new_n387), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n197), .A2(new_n198), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT83), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n197), .A2(KEYINPUT83), .A3(new_n198), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(KEYINPUT19), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT19), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n227), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n508), .A2(new_n204), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT82), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(new_n257), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n513), .B1(G214), .B2(new_n322), .ZN(new_n514));
  INV_X1    g328(.A(G237), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(new_n188), .A3(G214), .ZN(new_n516));
  NOR2_X1   g330(.A1(KEYINPUT82), .A2(G143), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(G131), .B1(new_n514), .B2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n516), .A2(new_n517), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n513), .A2(G214), .A3(new_n322), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(new_n521), .A3(new_n277), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n202), .A2(G146), .B1(new_n519), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n511), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g338(.A1(KEYINPUT18), .A2(G131), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n520), .A2(new_n521), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT84), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n520), .A2(new_n521), .A3(KEYINPUT84), .A4(new_n525), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n197), .A2(KEYINPUT83), .A3(new_n198), .ZN(new_n532));
  AOI21_X1  g346(.A(KEYINPUT83), .B1(new_n197), .B2(new_n198), .ZN(new_n533));
  NOR3_X1   g347(.A1(new_n532), .A2(new_n533), .A3(new_n204), .ZN(new_n534));
  INV_X1    g348(.A(new_n228), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n531), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n503), .B1(new_n524), .B2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT17), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n519), .A2(new_n538), .A3(new_n522), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n527), .A2(KEYINPUT17), .A3(G131), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n203), .A2(new_n539), .A3(new_n205), .A4(new_n540), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n536), .A2(new_n541), .A3(new_n503), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n501), .B1(new_n537), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(G475), .A2(G902), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n536), .A2(new_n541), .A3(new_n503), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n506), .A2(G146), .A3(new_n507), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n228), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n511), .A2(new_n523), .B1(new_n547), .B2(new_n531), .ZN(new_n548));
  OAI211_X1 g362(.A(KEYINPUT85), .B(new_n545), .C1(new_n548), .C2(new_n503), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n543), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT20), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT86), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n550), .A2(KEYINPUT86), .A3(KEYINPUT20), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n545), .B1(new_n548), .B2(new_n503), .ZN(new_n555));
  NOR3_X1   g369(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n553), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n503), .B1(new_n536), .B2(new_n541), .ZN(new_n559));
  AOI21_X1  g373(.A(G902), .B1(new_n559), .B2(KEYINPUT87), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n542), .A2(KEYINPUT87), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n560), .B1(new_n561), .B2(new_n559), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(G475), .ZN(new_n563));
  INV_X1    g377(.A(G478), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(KEYINPUT15), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT92), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n498), .A2(new_n240), .A3(G953), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT89), .B1(new_n218), .B2(G143), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT89), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(new_n257), .A3(G128), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n218), .A2(G143), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n571), .A2(new_n270), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT88), .B1(new_n310), .B2(G122), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT88), .ZN(new_n575));
  INV_X1    g389(.A(G122), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(G116), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n310), .A2(G122), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G107), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n390), .A3(new_n579), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n573), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT13), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n571), .A2(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n568), .A2(new_n570), .A3(KEYINPUT13), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n586), .A3(new_n572), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(G134), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n576), .A2(G116), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT14), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n590), .A2(KEYINPUT90), .A3(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(new_n310), .A3(G122), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT90), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n579), .A2(KEYINPUT14), .ZN(new_n596));
  NAND4_X1  g410(.A1(new_n578), .A2(new_n592), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(G107), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n270), .B1(new_n571), .B2(new_n572), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n598), .B(new_n582), .C1(new_n573), .C2(new_n599), .ZN(new_n600));
  AOI211_X1 g414(.A(new_n566), .B(new_n567), .C1(new_n589), .C2(new_n600), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n571), .A2(new_n584), .B1(new_n218), .B2(G143), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n270), .B1(new_n602), .B2(new_n586), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n571), .A2(new_n270), .A3(new_n572), .ZN(new_n604));
  AOI211_X1 g418(.A(G107), .B(new_n590), .C1(new_n577), .C2(new_n574), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n390), .B1(new_n578), .B2(new_n579), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n582), .B1(new_n573), .B2(new_n599), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n592), .A2(new_n595), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n574), .A2(new_n577), .B1(new_n579), .B2(KEYINPUT14), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n390), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  OAI22_X1  g425(.A1(new_n603), .A2(new_n607), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(new_n567), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT92), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n601), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n571), .A2(new_n572), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(G134), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n605), .B1(new_n617), .B2(new_n604), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n588), .A2(new_n583), .B1(new_n618), .B2(new_n598), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(KEYINPUT91), .A3(new_n567), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT91), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n621), .B1(new_n612), .B2(new_n613), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  AOI211_X1 g437(.A(G902), .B(new_n565), .C1(new_n615), .C2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(new_n565), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n566), .B1(new_n619), .B2(new_n567), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n567), .B1(new_n589), .B2(new_n600), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(KEYINPUT92), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT91), .B1(new_n619), .B2(new_n567), .ZN(new_n629));
  AND4_X1   g443(.A1(KEYINPUT91), .A2(new_n589), .A3(new_n600), .A4(new_n567), .ZN(new_n630));
  OAI211_X1 g444(.A(new_n626), .B(new_n628), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n625), .B1(new_n631), .B2(new_n241), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n624), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(G952), .ZN(new_n634));
  AOI211_X1 g448(.A(G953), .B(new_n634), .C1(G234), .C2(G237), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT21), .B(G898), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT93), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  AOI211_X1 g452(.A(new_n241), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n635), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n558), .A2(new_n563), .A3(new_n633), .A4(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n500), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n382), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n644), .B(G101), .ZN(G3));
  NAND2_X1  g459(.A1(new_n447), .A2(new_n499), .ZN(new_n646));
  INV_X1    g460(.A(G472), .ZN(new_n647));
  AOI21_X1  g461(.A(G902), .B1(new_n357), .B2(new_n358), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n250), .B(new_n349), .C1(new_n647), .C2(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(new_n650), .B(KEYINPUT94), .Z(new_n651));
  NOR2_X1   g465(.A1(new_n612), .A2(new_n613), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT33), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n652), .A2(new_n627), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n631), .B2(new_n653), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(G478), .A3(new_n241), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n631), .A2(new_n241), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n564), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n550), .A2(KEYINPUT86), .A3(KEYINPUT20), .ZN(new_n660));
  AOI21_X1  g474(.A(KEYINPUT86), .B1(new_n550), .B2(KEYINPUT20), .ZN(new_n661));
  INV_X1    g475(.A(new_n557), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n660), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(new_n563), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n659), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n448), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(new_n476), .B2(new_n487), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n496), .B1(new_n667), .B2(new_n493), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n641), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n651), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G104), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT95), .B(KEYINPUT34), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G6));
  INV_X1    g488(.A(KEYINPUT96), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n660), .B2(new_n661), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n553), .A2(KEYINPUT96), .A3(new_n554), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n543), .A2(new_n549), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n556), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n633), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n669), .A2(new_n664), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n651), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g498(.A(KEYINPUT35), .B(G107), .Z(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G9));
  NOR2_X1   g500(.A1(new_n648), .A2(new_n647), .ZN(new_n687));
  INV_X1    g501(.A(new_n242), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n688), .B1(new_n247), .B2(new_n248), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n236), .A2(new_n238), .ZN(new_n690));
  NOR2_X1   g504(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n692), .A2(new_n243), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n689), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n687), .A2(new_n694), .A3(new_n359), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n643), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT37), .B(G110), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G12));
  NAND2_X1  g512(.A1(new_n357), .A2(new_n358), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n360), .B1(new_n699), .B2(new_n252), .ZN(new_n700));
  AOI211_X1 g514(.A(KEYINPUT32), .B(new_n351), .C1(new_n357), .C2(new_n358), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n381), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n694), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n445), .B1(new_n432), .B2(new_n439), .ZN(new_n705));
  INV_X1    g519(.A(new_n499), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n668), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n704), .A2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT97), .ZN(new_n710));
  INV_X1    g524(.A(G900), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n635), .B1(new_n639), .B2(new_n711), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n712), .B1(new_n562), .B2(G475), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n680), .A2(new_n710), .A3(new_n681), .A4(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n680), .A2(new_n681), .A3(new_n713), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT97), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n709), .A2(new_n714), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G128), .ZN(G30));
  XOR2_X1   g532(.A(new_n712), .B(KEYINPUT39), .Z(new_n719));
  AND2_X1   g533(.A1(new_n707), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT40), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NOR3_X1   g536(.A1(new_n703), .A2(new_n633), .A3(new_n496), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n494), .B(KEYINPUT38), .Z(new_n724));
  NAND2_X1  g538(.A1(new_n558), .A2(new_n563), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n723), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n328), .A2(new_n334), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n356), .B1(new_n366), .B2(new_n367), .ZN(new_n729));
  AND2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(G472), .B1(new_n730), .B2(G902), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n362), .A2(KEYINPUT98), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT98), .B1(new_n362), .B2(new_n731), .ZN(new_n734));
  OR2_X1    g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n720), .A2(new_n721), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n727), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G143), .ZN(G45));
  INV_X1    g552(.A(new_n712), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n725), .A2(new_n659), .A3(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n709), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G146), .ZN(G48));
  INV_X1    g557(.A(KEYINPUT99), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n437), .A2(new_n241), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n744), .B1(new_n745), .B2(G469), .ZN(new_n746));
  AOI211_X1 g560(.A(KEYINPUT99), .B(new_n383), .C1(new_n437), .C2(new_n241), .ZN(new_n747));
  OAI211_X1 g561(.A(new_n440), .B(new_n499), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n382), .A2(new_n670), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT41), .B(G113), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n750), .B(new_n751), .ZN(G15));
  NAND3_X1  g566(.A1(new_n683), .A2(new_n382), .A3(new_n749), .ZN(new_n753));
  XOR2_X1   g567(.A(KEYINPUT100), .B(G116), .Z(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G18));
  INV_X1    g569(.A(KEYINPUT101), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n647), .B1(new_n376), .B2(new_n379), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n757), .B1(new_n350), .B2(new_n361), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n758), .A2(new_n642), .A3(new_n694), .ZN(new_n759));
  INV_X1    g573(.A(new_n668), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n748), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n756), .B1(new_n759), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n745), .A2(G469), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(KEYINPUT99), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n745), .A2(new_n744), .A3(G469), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(new_n499), .A3(new_n440), .A4(new_n668), .ZN(new_n767));
  NOR4_X1   g581(.A1(new_n704), .A2(new_n767), .A3(KEYINPUT101), .A4(new_n642), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n762), .A2(new_n768), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT102), .B(G119), .Z(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G21));
  NAND3_X1  g585(.A1(new_n364), .A2(new_n368), .A3(new_n372), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(new_n356), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT103), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n358), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n338), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n774), .B1(new_n773), .B2(new_n358), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n252), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n687), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n250), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n725), .A2(new_n681), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n640), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(new_n783), .A3(new_n761), .ZN(new_n784));
  XNOR2_X1  g598(.A(KEYINPUT104), .B(G122), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n784), .B(new_n785), .ZN(G24));
  NAND3_X1  g600(.A1(new_n778), .A2(new_n779), .A3(new_n703), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n787), .A2(new_n740), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n761), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G125), .ZN(G27));
  AND3_X1   g604(.A1(new_n488), .A2(new_n495), .A3(new_n493), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n702), .A2(new_n250), .A3(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n447), .A2(KEYINPUT105), .A3(new_n499), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT105), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n705), .B2(new_n706), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  AND4_X1   g610(.A1(KEYINPUT42), .A2(new_n792), .A3(new_n796), .A4(new_n741), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n702), .A2(new_n250), .A3(new_n791), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n793), .A2(new_n795), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT42), .B1(new_n801), .B2(new_n741), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G131), .ZN(G33));
  NAND4_X1  g619(.A1(new_n716), .A2(new_n792), .A3(new_n796), .A4(new_n714), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G134), .ZN(G36));
  OAI21_X1  g621(.A(new_n418), .B1(new_n435), .B2(new_n427), .ZN(new_n808));
  INV_X1    g622(.A(new_n386), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n808), .A2(new_n809), .B1(new_n441), .B2(new_n415), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT45), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(KEYINPUT45), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(G469), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(G469), .A2(G902), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT46), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n813), .A2(KEYINPUT46), .A3(new_n814), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n817), .A2(new_n440), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n499), .A3(new_n719), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n820), .A2(KEYINPUT106), .ZN(new_n821));
  INV_X1    g635(.A(new_n659), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n725), .A2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT43), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n694), .B1(new_n779), .B2(new_n349), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n824), .A2(KEYINPUT44), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n820), .A2(KEYINPUT106), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n821), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  AOI21_X1  g642(.A(KEYINPUT44), .B1(new_n824), .B2(new_n825), .ZN(new_n829));
  INV_X1    g643(.A(new_n791), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n828), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(G137), .ZN(G39));
  NOR4_X1   g647(.A1(new_n740), .A2(new_n702), .A3(new_n250), .A4(new_n830), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n819), .A2(KEYINPUT47), .A3(new_n499), .ZN(new_n835));
  AOI21_X1  g649(.A(KEYINPUT47), .B1(new_n819), .B2(new_n499), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n837), .B(G140), .ZN(G42));
  NAND4_X1  g652(.A1(new_n725), .A2(new_n681), .A3(new_n694), .A4(new_n739), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n839), .A2(new_n708), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n840), .B1(new_n733), .B2(new_n734), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n717), .A2(new_n841), .A3(new_n742), .A4(new_n789), .ZN(new_n842));
  XNOR2_X1  g656(.A(new_n842), .B(KEYINPUT52), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n844));
  INV_X1    g658(.A(new_n642), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n761), .A2(new_n845), .A3(new_n702), .A4(new_n703), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT101), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n382), .B(new_n749), .C1(new_n683), .C2(new_n670), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n848), .A2(new_n784), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n497), .A2(new_n641), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n646), .A2(new_n649), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT109), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n657), .A2(new_n565), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n631), .A2(new_n241), .A3(new_n625), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(KEYINPUT108), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT108), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n856), .B1(new_n624), .B2(new_n632), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n558), .A3(new_n563), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n852), .B1(new_n665), .B2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n859), .A2(new_n852), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n851), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n643), .B1(new_n382), .B2(new_n695), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n862), .A2(KEYINPUT110), .A3(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT110), .B1(new_n862), .B2(new_n863), .ZN(new_n865));
  OAI211_X1 g679(.A(new_n847), .B(new_n849), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n793), .A2(new_n795), .A3(new_n791), .ZN(new_n867));
  AND4_X1   g681(.A1(new_n713), .A2(new_n791), .A3(new_n855), .A4(new_n857), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n868), .A2(new_n680), .A3(new_n707), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n694), .B1(new_n362), .B2(new_n381), .ZN(new_n870));
  AOI22_X1  g684(.A1(new_n788), .A2(new_n867), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n806), .B(new_n871), .C1(new_n797), .C2(new_n802), .ZN(new_n872));
  NOR4_X1   g686(.A1(new_n843), .A2(new_n844), .A3(new_n866), .A4(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(new_n843), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n784), .B(new_n848), .C1(new_n762), .C2(new_n768), .ZN(new_n875));
  INV_X1    g689(.A(new_n865), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n862), .A2(new_n863), .A3(KEYINPUT110), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n871), .A2(new_n806), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n879), .B1(new_n803), .B2(new_n798), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT111), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT111), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n866), .A2(new_n882), .A3(new_n872), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n874), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT114), .ZN(new_n885));
  XNOR2_X1  g699(.A(KEYINPUT113), .B(KEYINPUT53), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  OAI21_X1  g701(.A(new_n882), .B1(new_n866), .B2(new_n872), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n876), .A2(new_n877), .ZN(new_n889));
  INV_X1    g703(.A(new_n875), .ZN(new_n890));
  NAND4_X1  g704(.A1(new_n880), .A2(new_n889), .A3(new_n890), .A4(KEYINPUT111), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n843), .B1(new_n888), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n886), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT114), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n873), .B1(new_n887), .B2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT54), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n888), .A2(new_n891), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n843), .B1(new_n898), .B2(KEYINPUT112), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(KEYINPUT112), .B2(new_n898), .ZN(new_n900));
  AOI22_X1  g714(.A1(new_n900), .A2(new_n844), .B1(new_n892), .B2(new_n893), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n897), .B1(new_n901), .B2(new_n896), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n824), .A2(new_n635), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n748), .A2(new_n830), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n905), .A2(new_n787), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n906), .B(KEYINPUT116), .Z(new_n907));
  AND2_X1   g721(.A1(new_n903), .A2(new_n781), .ZN(new_n908));
  INV_X1    g722(.A(new_n724), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT50), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n495), .B1(KEYINPUT115), .B2(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n908), .A2(new_n909), .A3(new_n749), .A4(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n910), .A2(KEYINPUT115), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n835), .A2(new_n836), .ZN(new_n915));
  AOI22_X1  g729(.A1(new_n764), .A2(new_n765), .B1(new_n439), .B2(new_n432), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n499), .B2(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n908), .A2(new_n791), .ZN(new_n919));
  AOI22_X1  g733(.A1(new_n918), .A2(new_n919), .B1(new_n912), .B2(new_n913), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n904), .A2(new_n250), .A3(new_n635), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n735), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n725), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n923), .A3(new_n822), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT117), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n907), .A2(new_n914), .A3(new_n920), .A4(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT51), .ZN(new_n927));
  OR2_X1    g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n908), .A2(new_n761), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT118), .ZN(new_n931));
  INV_X1    g745(.A(new_n382), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n905), .A2(new_n932), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT48), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n188), .A2(G952), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n735), .A2(new_n665), .A3(new_n921), .ZN(new_n936));
  NOR4_X1   g750(.A1(new_n931), .A2(new_n934), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n928), .A2(new_n929), .A3(new_n937), .ZN(new_n938));
  OAI22_X1  g752(.A1(new_n902), .A2(new_n938), .B1(G952), .B2(G953), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n659), .A2(new_n495), .A3(new_n499), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n724), .A2(new_n251), .A3(new_n940), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n917), .A2(KEYINPUT49), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n941), .A2(new_n923), .A3(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n917), .A2(KEYINPUT49), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n735), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT107), .Z(new_n946));
  NAND2_X1  g760(.A1(new_n939), .A2(new_n946), .ZN(G75));
  NOR2_X1   g761(.A1(new_n188), .A2(G952), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n948), .B(KEYINPUT121), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n895), .A2(new_n241), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n950), .A2(new_n449), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n474), .A2(new_n458), .A3(new_n475), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n492), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT55), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n954), .A2(KEYINPUT56), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n949), .B1(new_n951), .B2(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n873), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n885), .B1(new_n884), .B2(new_n886), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n892), .A2(KEYINPUT114), .A3(new_n893), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(G210), .A2(G902), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n960), .A2(KEYINPUT119), .A3(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT119), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n895), .B2(new_n961), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT56), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n963), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n954), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT120), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n967), .A2(KEYINPUT120), .A3(new_n954), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n956), .B1(new_n970), .B2(new_n971), .ZN(G51));
  NAND2_X1  g786(.A1(new_n960), .A2(KEYINPUT54), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n897), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n814), .B(KEYINPUT57), .Z(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n437), .ZN(new_n977));
  OR3_X1    g791(.A1(new_n895), .A2(new_n241), .A3(new_n813), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n948), .B1(new_n977), .B2(new_n978), .ZN(G54));
  AND2_X1   g793(.A1(KEYINPUT58), .A2(G475), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n950), .A2(new_n678), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n678), .B1(new_n950), .B2(new_n980), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n981), .A2(new_n982), .A3(new_n948), .ZN(G60));
  NAND2_X1  g797(.A1(G478), .A2(G902), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT59), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n974), .A2(new_n655), .A3(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n949), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n655), .B1(new_n902), .B2(new_n985), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(G63));
  NAND2_X1  g803(.A1(G217), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT122), .Z(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT60), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n895), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n692), .ZN(new_n994));
  INV_X1    g808(.A(new_n239), .ZN(new_n995));
  INV_X1    g809(.A(new_n233), .ZN(new_n996));
  OAI22_X1  g810(.A1(new_n895), .A2(new_n992), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n994), .A2(new_n949), .A3(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT61), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n998), .B(new_n999), .ZN(G66));
  OAI21_X1  g814(.A(G953), .B1(new_n638), .B2(new_n450), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n1001), .B1(new_n878), .B2(G953), .ZN(new_n1002));
  OAI211_X1 g816(.A(new_n474), .B(new_n475), .C1(G898), .C2(new_n188), .ZN(new_n1003));
  XNOR2_X1  g817(.A(new_n1002), .B(new_n1003), .ZN(G69));
  NOR3_X1   g818(.A1(new_n932), .A2(new_n760), .A3(new_n782), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n821), .A2(new_n827), .A3(new_n1005), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n1006), .A2(new_n806), .A3(new_n837), .ZN(new_n1007));
  AND3_X1   g821(.A1(new_n717), .A2(new_n742), .A3(new_n789), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1007), .A2(new_n832), .A3(new_n804), .A4(new_n1008), .ZN(new_n1009));
  OR2_X1    g823(.A1(new_n1009), .A2(KEYINPUT125), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(KEYINPUT125), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n1010), .A2(new_n188), .A3(new_n1011), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n298), .A2(new_n308), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n508), .A2(new_n510), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(G900), .A2(G953), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1012), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT124), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1008), .A2(new_n737), .ZN(new_n1019));
  OR2_X1    g833(.A1(new_n1019), .A2(KEYINPUT62), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n792), .B(new_n720), .C1(new_n860), .C2(new_n861), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n837), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n1022), .B1(new_n828), .B2(new_n831), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1019), .A2(KEYINPUT62), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1020), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT123), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n1020), .A2(new_n1023), .A3(KEYINPUT123), .A4(new_n1024), .ZN(new_n1028));
  AOI21_X1  g842(.A(G953), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1018), .B1(new_n1029), .B2(new_n1015), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1017), .A2(new_n1030), .ZN(new_n1031));
  NOR3_X1   g845(.A1(new_n1029), .A2(new_n1018), .A3(new_n1015), .ZN(new_n1032));
  OAI21_X1  g846(.A(KEYINPUT126), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1032), .ZN(new_n1035));
  INV_X1    g849(.A(KEYINPUT126), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n1035), .A2(new_n1036), .A3(new_n1017), .A4(new_n1030), .ZN(new_n1037));
  AND3_X1   g851(.A1(new_n1033), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1034), .B1(new_n1033), .B2(new_n1037), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1038), .A2(new_n1039), .ZN(G72));
  NAND2_X1  g854(.A1(G472), .A2(G902), .ZN(new_n1041));
  XOR2_X1   g855(.A(new_n1041), .B(KEYINPUT63), .Z(new_n1042));
  INV_X1    g856(.A(new_n1042), .ZN(new_n1043));
  AOI211_X1 g857(.A(new_n1043), .B(new_n901), .C1(new_n728), .C2(new_n378), .ZN(new_n1044));
  INV_X1    g858(.A(new_n377), .ZN(new_n1045));
  NAND3_X1  g859(.A1(new_n1027), .A2(new_n878), .A3(new_n1028), .ZN(new_n1046));
  AOI211_X1 g860(.A(new_n356), .B(new_n1045), .C1(new_n1046), .C2(new_n1042), .ZN(new_n1047));
  XNOR2_X1  g861(.A(new_n1047), .B(KEYINPUT127), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1010), .A2(new_n878), .A3(new_n1011), .ZN(new_n1049));
  AOI211_X1 g863(.A(new_n326), .B(new_n377), .C1(new_n1049), .C2(new_n1042), .ZN(new_n1050));
  NOR4_X1   g864(.A1(new_n1044), .A2(new_n1048), .A3(new_n948), .A4(new_n1050), .ZN(G57));
endmodule


