

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585;

  OR2_X1 U320 ( .A1(n442), .A2(n445), .ZN(n444) );
  XNOR2_X1 U321 ( .A(n314), .B(n313), .ZN(n315) );
  NOR2_X1 U322 ( .A1(n474), .A2(n501), .ZN(n567) );
  XOR2_X1 U323 ( .A(KEYINPUT26), .B(n423), .Z(n565) );
  XNOR2_X1 U324 ( .A(n458), .B(KEYINPUT64), .ZN(n459) );
  XNOR2_X1 U325 ( .A(n460), .B(n459), .ZN(n461) );
  INV_X1 U326 ( .A(G190GAT), .ZN(n370) );
  XNOR2_X1 U327 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U328 ( .A(n437), .B(n372), .ZN(n373) );
  INV_X1 U329 ( .A(KEYINPUT72), .ZN(n311) );
  INV_X1 U330 ( .A(KEYINPUT99), .ZN(n443) );
  XNOR2_X1 U331 ( .A(n312), .B(n311), .ZN(n313) );
  NOR2_X1 U332 ( .A1(n385), .A2(n475), .ZN(n423) );
  XNOR2_X1 U333 ( .A(KEYINPUT102), .B(KEYINPUT36), .ZN(n361) );
  XNOR2_X1 U334 ( .A(n357), .B(n356), .ZN(n358) );
  NOR2_X1 U335 ( .A1(n562), .A2(n450), .ZN(n451) );
  XNOR2_X1 U336 ( .A(n483), .B(n361), .ZN(n581) );
  XNOR2_X1 U337 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U338 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U339 ( .A(n321), .B(n320), .ZN(n572) );
  XNOR2_X1 U340 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U341 ( .A(n455), .B(G43GAT), .ZN(n456) );
  XNOR2_X1 U342 ( .A(n487), .B(n486), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(n457), .B(n456), .ZN(G1330GAT) );
  XOR2_X1 U344 ( .A(KEYINPUT38), .B(KEYINPUT103), .Z(n453) );
  XOR2_X1 U345 ( .A(G169GAT), .B(G8GAT), .Z(n391) );
  XOR2_X1 U346 ( .A(G141GAT), .B(G50GAT), .Z(n289) );
  XNOR2_X1 U347 ( .A(G36GAT), .B(G29GAT), .ZN(n288) );
  XNOR2_X1 U348 ( .A(n289), .B(n288), .ZN(n290) );
  XOR2_X1 U349 ( .A(n391), .B(n290), .Z(n292) );
  NAND2_X1 U350 ( .A1(G229GAT), .A2(G233GAT), .ZN(n291) );
  XNOR2_X1 U351 ( .A(n292), .B(n291), .ZN(n305) );
  XOR2_X1 U352 ( .A(G197GAT), .B(KEYINPUT67), .Z(n294) );
  XNOR2_X1 U353 ( .A(KEYINPUT65), .B(KEYINPUT69), .ZN(n293) );
  XNOR2_X1 U354 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U355 ( .A(KEYINPUT30), .B(KEYINPUT66), .Z(n296) );
  XNOR2_X1 U356 ( .A(G113GAT), .B(KEYINPUT29), .ZN(n295) );
  XNOR2_X1 U357 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U358 ( .A(n298), .B(n297), .Z(n303) );
  XNOR2_X1 U359 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n299) );
  XNOR2_X1 U360 ( .A(n299), .B(KEYINPUT7), .ZN(n355) );
  XOR2_X1 U361 ( .A(G1GAT), .B(G15GAT), .Z(n301) );
  XNOR2_X1 U362 ( .A(KEYINPUT68), .B(G22GAT), .ZN(n300) );
  XNOR2_X1 U363 ( .A(n301), .B(n300), .ZN(n331) );
  XNOR2_X1 U364 ( .A(n355), .B(n331), .ZN(n302) );
  XNOR2_X1 U365 ( .A(n303), .B(n302), .ZN(n304) );
  XNOR2_X1 U366 ( .A(n305), .B(n304), .ZN(n568) );
  INV_X1 U367 ( .A(n568), .ZN(n560) );
  XNOR2_X1 U368 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n306) );
  XNOR2_X1 U369 ( .A(n306), .B(G78GAT), .ZN(n329) );
  XOR2_X1 U370 ( .A(G99GAT), .B(G106GAT), .Z(n356) );
  XOR2_X1 U371 ( .A(n329), .B(n356), .Z(n308) );
  NAND2_X1 U372 ( .A1(G230GAT), .A2(G233GAT), .ZN(n307) );
  XNOR2_X1 U373 ( .A(n308), .B(n307), .ZN(n314) );
  XOR2_X1 U374 ( .A(G64GAT), .B(G204GAT), .Z(n310) );
  XNOR2_X1 U375 ( .A(G176GAT), .B(KEYINPUT71), .ZN(n309) );
  XNOR2_X1 U376 ( .A(n310), .B(n309), .ZN(n397) );
  XNOR2_X1 U377 ( .A(n397), .B(KEYINPUT31), .ZN(n312) );
  XOR2_X1 U378 ( .A(G120GAT), .B(G57GAT), .Z(n431) );
  XOR2_X1 U379 ( .A(n315), .B(n431), .Z(n321) );
  XOR2_X1 U380 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n317) );
  XNOR2_X1 U381 ( .A(G148GAT), .B(KEYINPUT70), .ZN(n316) );
  XOR2_X1 U382 ( .A(n317), .B(n316), .Z(n319) );
  XNOR2_X1 U383 ( .A(G92GAT), .B(G85GAT), .ZN(n318) );
  AND2_X1 U384 ( .A1(n560), .A2(n572), .ZN(n491) );
  XOR2_X1 U385 ( .A(KEYINPUT77), .B(KEYINPUT14), .Z(n323) );
  XNOR2_X1 U386 ( .A(KEYINPUT15), .B(KEYINPUT12), .ZN(n322) );
  XNOR2_X1 U387 ( .A(n323), .B(n322), .ZN(n339) );
  XOR2_X1 U388 ( .A(KEYINPUT80), .B(KEYINPUT78), .Z(n325) );
  XNOR2_X1 U389 ( .A(G8GAT), .B(KEYINPUT79), .ZN(n324) );
  XNOR2_X1 U390 ( .A(n325), .B(n324), .ZN(n327) );
  XOR2_X1 U391 ( .A(G57GAT), .B(G64GAT), .Z(n326) );
  XNOR2_X1 U392 ( .A(n327), .B(n326), .ZN(n335) );
  XNOR2_X1 U393 ( .A(G127GAT), .B(G211GAT), .ZN(n328) );
  XNOR2_X1 U394 ( .A(n328), .B(G155GAT), .ZN(n330) );
  XOR2_X1 U395 ( .A(n330), .B(n329), .Z(n333) );
  XNOR2_X1 U396 ( .A(n331), .B(G183GAT), .ZN(n332) );
  XNOR2_X1 U397 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U398 ( .A(n335), .B(n334), .ZN(n337) );
  NAND2_X1 U399 ( .A1(G231GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U400 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U401 ( .A(n339), .B(n338), .ZN(n562) );
  XOR2_X1 U402 ( .A(G218GAT), .B(G92GAT), .Z(n341) );
  XNOR2_X1 U403 ( .A(G36GAT), .B(G190GAT), .ZN(n340) );
  XNOR2_X1 U404 ( .A(n341), .B(n340), .ZN(n387) );
  INV_X1 U405 ( .A(KEYINPUT74), .ZN(n342) );
  XNOR2_X1 U406 ( .A(n387), .B(n342), .ZN(n346) );
  INV_X1 U407 ( .A(n346), .ZN(n344) );
  NAND2_X1 U408 ( .A1(G232GAT), .A2(G233GAT), .ZN(n345) );
  INV_X1 U409 ( .A(n345), .ZN(n343) );
  NAND2_X1 U410 ( .A1(n344), .A2(n343), .ZN(n348) );
  NAND2_X1 U411 ( .A1(n346), .A2(n345), .ZN(n347) );
  NAND2_X1 U412 ( .A1(n348), .A2(n347), .ZN(n352) );
  XOR2_X1 U413 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n350) );
  XNOR2_X1 U414 ( .A(KEYINPUT11), .B(KEYINPUT73), .ZN(n349) );
  XOR2_X1 U415 ( .A(n350), .B(n349), .Z(n351) );
  XNOR2_X1 U416 ( .A(n352), .B(n351), .ZN(n359) );
  XOR2_X1 U417 ( .A(KEYINPUT75), .B(G85GAT), .Z(n354) );
  XNOR2_X1 U418 ( .A(G29GAT), .B(G134GAT), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n354), .B(n353), .ZN(n436) );
  XNOR2_X1 U420 ( .A(n355), .B(n436), .ZN(n357) );
  XNOR2_X1 U421 ( .A(G50GAT), .B(G162GAT), .ZN(n405) );
  XNOR2_X1 U422 ( .A(n360), .B(n405), .ZN(n557) );
  XNOR2_X1 U423 ( .A(KEYINPUT76), .B(n557), .ZN(n483) );
  XOR2_X1 U424 ( .A(G120GAT), .B(G71GAT), .Z(n363) );
  XNOR2_X1 U425 ( .A(G169GAT), .B(G176GAT), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U427 ( .A(KEYINPUT84), .B(KEYINPUT86), .Z(n365) );
  XNOR2_X1 U428 ( .A(G15GAT), .B(KEYINPUT87), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U430 ( .A(n367), .B(n366), .Z(n375) );
  XOR2_X1 U431 ( .A(KEYINPUT0), .B(KEYINPUT81), .Z(n369) );
  XNOR2_X1 U432 ( .A(G113GAT), .B(G127GAT), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n369), .B(n368), .ZN(n437) );
  XNOR2_X1 U434 ( .A(G43GAT), .B(G134GAT), .ZN(n371) );
  XNOR2_X1 U435 ( .A(G99GAT), .B(n373), .ZN(n374) );
  XNOR2_X1 U436 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U437 ( .A(KEYINPUT83), .B(KEYINPUT82), .Z(n377) );
  NAND2_X1 U438 ( .A1(G227GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U440 ( .A(n379), .B(n378), .Z(n384) );
  XOR2_X1 U441 ( .A(KEYINPUT17), .B(G183GAT), .Z(n381) );
  XNOR2_X1 U442 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U444 ( .A(KEYINPUT85), .B(n382), .Z(n398) );
  XNOR2_X1 U445 ( .A(n398), .B(KEYINPUT20), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n384), .B(n383), .ZN(n385) );
  INV_X1 U447 ( .A(n385), .ZN(n386) );
  XOR2_X1 U448 ( .A(n387), .B(KEYINPUT97), .Z(n389) );
  NAND2_X1 U449 ( .A1(G226GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U450 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U451 ( .A(n390), .B(KEYINPUT96), .Z(n393) );
  XNOR2_X1 U452 ( .A(n391), .B(KEYINPUT95), .ZN(n392) );
  XNOR2_X1 U453 ( .A(n393), .B(n392), .ZN(n396) );
  XOR2_X1 U454 ( .A(KEYINPUT91), .B(KEYINPUT21), .Z(n395) );
  XNOR2_X1 U455 ( .A(G197GAT), .B(G211GAT), .ZN(n394) );
  XNOR2_X1 U456 ( .A(n395), .B(n394), .ZN(n408) );
  XOR2_X1 U457 ( .A(n396), .B(n408), .Z(n400) );
  XNOR2_X1 U458 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U459 ( .A(n400), .B(n399), .ZN(n504) );
  NAND2_X1 U460 ( .A1(n385), .A2(n504), .ZN(n401) );
  XNOR2_X1 U461 ( .A(KEYINPUT98), .B(n401), .ZN(n421) );
  XOR2_X1 U462 ( .A(G218GAT), .B(G78GAT), .Z(n403) );
  XNOR2_X1 U463 ( .A(G204GAT), .B(G106GAT), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U465 ( .A(n404), .B(KEYINPUT90), .Z(n407) );
  XOR2_X1 U466 ( .A(G22GAT), .B(n405), .Z(n406) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n412) );
  XOR2_X1 U468 ( .A(n408), .B(KEYINPUT89), .Z(n410) );
  NAND2_X1 U469 ( .A1(G228GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U470 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U471 ( .A(n412), .B(n411), .Z(n420) );
  XOR2_X1 U472 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n414) );
  XNOR2_X1 U473 ( .A(G141GAT), .B(G148GAT), .ZN(n413) );
  XNOR2_X1 U474 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U475 ( .A(G155GAT), .B(n415), .Z(n434) );
  XOR2_X1 U476 ( .A(KEYINPUT22), .B(KEYINPUT88), .Z(n417) );
  XNOR2_X1 U477 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n416) );
  XNOR2_X1 U478 ( .A(n417), .B(n416), .ZN(n418) );
  XNOR2_X1 U479 ( .A(n434), .B(n418), .ZN(n419) );
  XNOR2_X1 U480 ( .A(n420), .B(n419), .ZN(n475) );
  NAND2_X1 U481 ( .A1(n421), .A2(n475), .ZN(n422) );
  XNOR2_X1 U482 ( .A(n422), .B(KEYINPUT25), .ZN(n425) );
  INV_X1 U483 ( .A(n504), .ZN(n522) );
  XNOR2_X1 U484 ( .A(n522), .B(KEYINPUT27), .ZN(n446) );
  NOR2_X1 U485 ( .A1(n446), .A2(n565), .ZN(n424) );
  NOR2_X1 U486 ( .A1(n425), .A2(n424), .ZN(n442) );
  XOR2_X1 U487 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n427) );
  XNOR2_X1 U488 ( .A(KEYINPUT93), .B(KEYINPUT4), .ZN(n426) );
  XNOR2_X1 U489 ( .A(n427), .B(n426), .ZN(n441) );
  XOR2_X1 U490 ( .A(KEYINPUT92), .B(KEYINPUT6), .Z(n429) );
  XNOR2_X1 U491 ( .A(G1GAT), .B(G162GAT), .ZN(n428) );
  XNOR2_X1 U492 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U493 ( .A(n431), .B(n430), .Z(n433) );
  NAND2_X1 U494 ( .A1(G225GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U495 ( .A(n433), .B(n432), .ZN(n435) );
  XOR2_X1 U496 ( .A(n435), .B(n434), .Z(n439) );
  XNOR2_X1 U497 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U499 ( .A(n441), .B(n440), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n449) );
  XOR2_X1 U501 ( .A(KEYINPUT94), .B(n445), .Z(n520) );
  NOR2_X1 U502 ( .A1(n446), .A2(n520), .ZN(n532) );
  XNOR2_X1 U503 ( .A(n475), .B(KEYINPUT28), .ZN(n527) );
  INV_X1 U504 ( .A(n527), .ZN(n534) );
  NOR2_X1 U505 ( .A1(n385), .A2(n534), .ZN(n447) );
  NAND2_X1 U506 ( .A1(n532), .A2(n447), .ZN(n448) );
  NAND2_X1 U507 ( .A1(n449), .A2(n448), .ZN(n489) );
  NAND2_X1 U508 ( .A1(n581), .A2(n489), .ZN(n450) );
  XOR2_X1 U509 ( .A(KEYINPUT37), .B(n451), .Z(n519) );
  NAND2_X1 U510 ( .A1(n491), .A2(n519), .ZN(n452) );
  XNOR2_X1 U511 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U512 ( .A(KEYINPUT104), .B(n454), .Z(n506) );
  NAND2_X1 U513 ( .A1(n506), .A2(n385), .ZN(n457) );
  XOR2_X1 U514 ( .A(KEYINPUT40), .B(KEYINPUT105), .Z(n455) );
  NAND2_X1 U515 ( .A1(n581), .A2(n562), .ZN(n460) );
  XOR2_X1 U516 ( .A(KEYINPUT45), .B(KEYINPUT110), .Z(n458) );
  NAND2_X1 U517 ( .A1(n461), .A2(n572), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT111), .ZN(n463) );
  NAND2_X1 U519 ( .A1(n463), .A2(n568), .ZN(n470) );
  INV_X1 U520 ( .A(n562), .ZN(n577) );
  XOR2_X1 U521 ( .A(KEYINPUT41), .B(n572), .Z(n508) );
  NOR2_X1 U522 ( .A1(n508), .A2(n568), .ZN(n465) );
  XNOR2_X1 U523 ( .A(KEYINPUT46), .B(KEYINPUT109), .ZN(n464) );
  XNOR2_X1 U524 ( .A(n465), .B(n464), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n577), .A2(n466), .ZN(n467) );
  NOR2_X1 U526 ( .A1(n557), .A2(n467), .ZN(n468) );
  XNOR2_X1 U527 ( .A(KEYINPUT47), .B(n468), .ZN(n469) );
  NAND2_X1 U528 ( .A1(n470), .A2(n469), .ZN(n471) );
  XNOR2_X1 U529 ( .A(n471), .B(KEYINPUT48), .ZN(n531) );
  XNOR2_X1 U530 ( .A(KEYINPUT119), .B(n522), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n531), .A2(n472), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n473), .B(KEYINPUT54), .ZN(n474) );
  INV_X1 U533 ( .A(n520), .ZN(n501) );
  NAND2_X1 U534 ( .A1(n567), .A2(n475), .ZN(n476) );
  XNOR2_X1 U535 ( .A(n476), .B(KEYINPUT55), .ZN(n477) );
  NAND2_X1 U536 ( .A1(n477), .A2(n385), .ZN(n478) );
  XOR2_X1 U537 ( .A(KEYINPUT120), .B(n478), .Z(n563) );
  INV_X1 U538 ( .A(n508), .ZN(n552) );
  NAND2_X1 U539 ( .A1(n563), .A2(n552), .ZN(n482) );
  XOR2_X1 U540 ( .A(G176GAT), .B(KEYINPUT121), .Z(n480) );
  XOR2_X1 U541 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n479) );
  XNOR2_X1 U542 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U543 ( .A(n482), .B(n481), .ZN(G1349GAT) );
  NAND2_X1 U544 ( .A1(n563), .A2(n483), .ZN(n487) );
  XOR2_X1 U545 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n485) );
  XNOR2_X1 U546 ( .A(G190GAT), .B(KEYINPUT122), .ZN(n484) );
  NOR2_X1 U547 ( .A1(n483), .A2(n577), .ZN(n488) );
  XNOR2_X1 U548 ( .A(KEYINPUT16), .B(n488), .ZN(n490) );
  AND2_X1 U549 ( .A1(n490), .A2(n489), .ZN(n509) );
  NAND2_X1 U550 ( .A1(n491), .A2(n509), .ZN(n499) );
  NOR2_X1 U551 ( .A1(n520), .A2(n499), .ZN(n492) );
  XOR2_X1 U552 ( .A(KEYINPUT34), .B(n492), .Z(n493) );
  XNOR2_X1 U553 ( .A(G1GAT), .B(n493), .ZN(G1324GAT) );
  NOR2_X1 U554 ( .A1(n522), .A2(n499), .ZN(n494) );
  XOR2_X1 U555 ( .A(G8GAT), .B(n494), .Z(G1325GAT) );
  NOR2_X1 U556 ( .A1(n499), .A2(n386), .ZN(n498) );
  XOR2_X1 U557 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n496) );
  XNOR2_X1 U558 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n495) );
  XNOR2_X1 U559 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1326GAT) );
  NOR2_X1 U561 ( .A1(n527), .A2(n499), .ZN(n500) );
  XOR2_X1 U562 ( .A(G22GAT), .B(n500), .Z(G1327GAT) );
  XOR2_X1 U563 ( .A(G29GAT), .B(KEYINPUT39), .Z(n503) );
  NAND2_X1 U564 ( .A1(n506), .A2(n501), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n503), .B(n502), .ZN(G1328GAT) );
  NAND2_X1 U566 ( .A1(n506), .A2(n504), .ZN(n505) );
  XNOR2_X1 U567 ( .A(n505), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U568 ( .A1(n506), .A2(n534), .ZN(n507) );
  XNOR2_X1 U569 ( .A(n507), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U570 ( .A1(n560), .A2(n508), .ZN(n518) );
  NAND2_X1 U571 ( .A1(n518), .A2(n509), .ZN(n515) );
  NOR2_X1 U572 ( .A1(n520), .A2(n515), .ZN(n510) );
  XOR2_X1 U573 ( .A(G57GAT), .B(n510), .Z(n511) );
  XNOR2_X1 U574 ( .A(KEYINPUT42), .B(n511), .ZN(G1332GAT) );
  NOR2_X1 U575 ( .A1(n522), .A2(n515), .ZN(n512) );
  XOR2_X1 U576 ( .A(G64GAT), .B(n512), .Z(G1333GAT) );
  NOR2_X1 U577 ( .A1(n386), .A2(n515), .ZN(n513) );
  XOR2_X1 U578 ( .A(KEYINPUT106), .B(n513), .Z(n514) );
  XNOR2_X1 U579 ( .A(G71GAT), .B(n514), .ZN(G1334GAT) );
  NOR2_X1 U580 ( .A1(n527), .A2(n515), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n526) );
  NOR2_X1 U584 ( .A1(n520), .A2(n526), .ZN(n521) );
  XOR2_X1 U585 ( .A(G85GAT), .B(n521), .Z(G1336GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n526), .ZN(n523) );
  XOR2_X1 U587 ( .A(G92GAT), .B(n523), .Z(G1337GAT) );
  NOR2_X1 U588 ( .A1(n386), .A2(n526), .ZN(n525) );
  XNOR2_X1 U589 ( .A(G99GAT), .B(KEYINPUT107), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1338GAT) );
  NOR2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U592 ( .A(KEYINPUT108), .B(KEYINPUT44), .ZN(n528) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(n530) );
  XOR2_X1 U594 ( .A(G106GAT), .B(n530), .Z(G1339GAT) );
  NAND2_X1 U595 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U596 ( .A(n533), .B(KEYINPUT112), .ZN(n549) );
  NOR2_X1 U597 ( .A1(n549), .A2(n534), .ZN(n535) );
  NAND2_X1 U598 ( .A1(n385), .A2(n535), .ZN(n536) );
  XNOR2_X1 U599 ( .A(KEYINPUT113), .B(n536), .ZN(n546) );
  NAND2_X1 U600 ( .A1(n546), .A2(n560), .ZN(n539) );
  XOR2_X1 U601 ( .A(G113GAT), .B(KEYINPUT114), .Z(n537) );
  XNOR2_X1 U602 ( .A(KEYINPUT115), .B(n537), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n541) );
  NAND2_X1 U605 ( .A1(n546), .A2(n552), .ZN(n540) );
  XNOR2_X1 U606 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(G120GAT), .B(n542), .ZN(G1341GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n544) );
  NAND2_X1 U609 ( .A1(n546), .A2(n562), .ZN(n543) );
  XNOR2_X1 U610 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U613 ( .A1(n546), .A2(n483), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1343GAT) );
  NOR2_X1 U615 ( .A1(n549), .A2(n565), .ZN(n550) );
  XNOR2_X1 U616 ( .A(KEYINPUT118), .B(n550), .ZN(n558) );
  NAND2_X1 U617 ( .A1(n558), .A2(n560), .ZN(n551) );
  XNOR2_X1 U618 ( .A(n551), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  NAND2_X1 U620 ( .A1(n558), .A2(n552), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n562), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U627 ( .A1(n560), .A2(n563), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G169GAT), .B(n561), .ZN(G1348GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G183GAT), .ZN(G1350GAT) );
  INV_X1 U631 ( .A(n565), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n580) );
  NOR2_X1 U633 ( .A1(n568), .A2(n580), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U637 ( .A1(n580), .A2(n572), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n574) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n580), .ZN(n578) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(n578), .Z(n579) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  XOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n584) );
  INV_X1 U646 ( .A(n580), .ZN(n582) );
  NAND2_X1 U647 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U648 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(n585), .ZN(G1355GAT) );
endmodule

