//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 0 0 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1253, new_n1254, new_n1255, new_n1256;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  AND2_X1   g0009(.A1(G116), .A2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G77), .ZN(new_n211));
  INV_X1    g0011(.A(G244), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI22_X1  g0014(.A1(new_n211), .A2(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n210), .B(new_n215), .C1(G87), .C2(G250), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G58), .A2(G232), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G107), .A2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G50), .A2(G226), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G68), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n209), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n209), .A2(G13), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n226), .B(G250), .C1(G257), .C2(G264), .ZN(new_n227));
  XOR2_X1   g0027(.A(new_n227), .B(KEYINPUT0), .Z(new_n228));
  OAI21_X1  g0028(.A(G50), .B1(G58), .B2(G68), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n229), .A2(new_n207), .A3(new_n230), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n225), .A2(new_n228), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT64), .ZN(new_n237));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(G264), .B(G270), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT65), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  AND2_X1   g0050(.A1(KEYINPUT3), .A2(G33), .ZN(new_n251));
  NOR2_X1   g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  OAI211_X1 g0052(.A(G226), .B(new_n250), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT69), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  OR2_X1    g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g0058(.A1(new_n258), .A2(KEYINPUT69), .A3(G226), .A4(new_n250), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G97), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n251), .A2(new_n252), .ZN(new_n262));
  INV_X1    g0062(.A(G232), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G1698), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n260), .A2(new_n261), .A3(new_n265), .ZN(new_n266));
  AND2_X1   g0066(.A1(G33), .A2(G41), .ZN(new_n267));
  OR2_X1    g0067(.A1(new_n267), .A2(new_n230), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n266), .A2(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  OR2_X1    g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n268), .A2(new_n271), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G238), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n270), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT13), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT13), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n270), .A2(new_n279), .A3(new_n273), .A4(new_n276), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n278), .A2(new_n280), .A3(KEYINPUT70), .ZN(new_n281));
  OR3_X1    g0081(.A1(new_n277), .A2(KEYINPUT70), .A3(KEYINPUT13), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n281), .A2(new_n282), .A3(G169), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(KEYINPUT14), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT14), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n281), .A2(new_n282), .A3(new_n285), .A4(G169), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n278), .A2(new_n280), .A3(G179), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n230), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(new_n206), .B2(G20), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT12), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n293), .B1(new_n295), .B2(new_n221), .ZN(new_n296));
  NOR3_X1   g0096(.A1(new_n294), .A2(KEYINPUT12), .A3(G68), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n292), .A2(new_n221), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT66), .ZN(new_n299));
  INV_X1    g0099(.A(G33), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n299), .A2(new_n207), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g0101(.A(KEYINPUT66), .B1(G20), .B2(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(G50), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT71), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n304), .B(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n207), .A2(G33), .ZN(new_n307));
  OAI221_X1 g0107(.A(new_n306), .B1(new_n207), .B2(G68), .C1(new_n211), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n290), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(KEYINPUT11), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT11), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n308), .A2(new_n311), .A3(new_n290), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n298), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n288), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n281), .A2(new_n282), .A3(G200), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n278), .A2(new_n280), .A3(G190), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n316), .A2(new_n313), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(KEYINPUT72), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT72), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n316), .A2(new_n313), .A3(new_n320), .A4(new_n317), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n294), .A2(G77), .ZN(new_n322));
  INV_X1    g0122(.A(new_n290), .ZN(new_n323));
  XOR2_X1   g0123(.A(KEYINPUT15), .B(G87), .Z(new_n324));
  INV_X1    g0124(.A(new_n307), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n324), .A2(new_n325), .B1(G20), .B2(G77), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT8), .B(G58), .Z(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n303), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n323), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  AOI211_X1 g0129(.A(new_n322), .B(new_n329), .C1(G77), .C2(new_n291), .ZN(new_n330));
  INV_X1    g0130(.A(new_n273), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n264), .A2(new_n250), .ZN(new_n332));
  INV_X1    g0132(.A(G107), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n250), .B1(new_n256), .B2(new_n257), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  OAI221_X1 g0135(.A(new_n332), .B1(new_n333), .B2(new_n258), .C1(new_n335), .C2(new_n222), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n331), .B1(new_n336), .B2(new_n269), .ZN(new_n337));
  INV_X1    g0137(.A(G179), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n275), .A2(G244), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT68), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n340), .A2(new_n341), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n330), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n337), .A2(new_n339), .ZN(new_n345));
  INV_X1    g0145(.A(G169), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n344), .A2(new_n347), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n315), .A2(new_n319), .A3(new_n321), .A4(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n327), .A2(new_n325), .B1(G20), .B2(new_n203), .ZN(new_n350));
  INV_X1    g0150(.A(G150), .ZN(new_n351));
  INV_X1    g0151(.A(new_n303), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n350), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n353), .A2(new_n290), .B1(new_n202), .B2(new_n295), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n202), .B2(new_n292), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT9), .ZN(new_n356));
  NOR2_X1   g0156(.A1(G222), .A2(G1698), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n250), .A2(G223), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n258), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(new_n269), .C1(G77), .C2(new_n258), .ZN(new_n360));
  INV_X1    g0160(.A(G226), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n360), .B(new_n273), .C1(new_n361), .C2(new_n274), .ZN(new_n362));
  XOR2_X1   g0162(.A(KEYINPUT67), .B(G200), .Z(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G190), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n356), .B(new_n364), .C1(new_n365), .C2(new_n362), .ZN(new_n366));
  XNOR2_X1  g0166(.A(new_n366), .B(KEYINPUT10), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n362), .A2(new_n346), .ZN(new_n368));
  OAI211_X1 g0168(.A(new_n355), .B(new_n368), .C1(G179), .C2(new_n362), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT18), .ZN(new_n371));
  INV_X1    g0171(.A(G87), .ZN(new_n372));
  NOR2_X1   g0172(.A1(new_n300), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(G223), .A2(G1698), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n374), .B1(new_n256), .B2(new_n257), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n361), .A2(G1698), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n373), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n377), .A2(new_n268), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT76), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n268), .A2(G232), .A3(new_n271), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .A4(new_n273), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(new_n273), .C1(new_n377), .C2(new_n268), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT76), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n381), .A2(new_n383), .A3(new_n346), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n382), .A2(G179), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g0186(.A(KEYINPUT8), .B(G58), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n294), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n388), .B1(new_n291), .B2(new_n387), .ZN(new_n389));
  XOR2_X1   g0189(.A(new_n389), .B(KEYINPUT75), .Z(new_n390));
  INV_X1    g0190(.A(KEYINPUT73), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n391), .B1(new_n303), .B2(G159), .ZN(new_n392));
  INV_X1    g0192(.A(G159), .ZN(new_n393));
  AOI211_X1 g0193(.A(KEYINPUT73), .B(new_n393), .C1(new_n301), .C2(new_n302), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT7), .B1(new_n262), .B2(new_n207), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NOR4_X1   g0197(.A1(new_n251), .A2(new_n252), .A3(new_n397), .A4(G20), .ZN(new_n398));
  OAI21_X1  g0198(.A(G68), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G58), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n400), .A2(new_n221), .ZN(new_n401));
  OAI21_X1  g0201(.A(G20), .B1(new_n401), .B2(new_n201), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n395), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n395), .A2(new_n399), .A3(KEYINPUT16), .A4(new_n402), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n405), .A2(new_n290), .A3(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT74), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n390), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n405), .A2(KEYINPUT74), .A3(new_n290), .A4(new_n406), .ZN(new_n410));
  AOI211_X1 g0210(.A(new_n371), .B(new_n386), .C1(new_n409), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n408), .ZN(new_n412));
  INV_X1    g0212(.A(new_n390), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n412), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n386), .ZN(new_n415));
  AOI21_X1  g0215(.A(KEYINPUT18), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G200), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n381), .A2(new_n383), .A3(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(G190), .B2(new_n382), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n409), .A2(new_n420), .A3(new_n410), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT17), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n409), .A2(new_n420), .A3(KEYINPUT17), .A4(new_n410), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OR2_X1    g0225(.A1(new_n417), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n345), .A2(new_n363), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n427), .B(new_n330), .C1(new_n365), .C2(new_n345), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NOR4_X1   g0229(.A1(new_n349), .A2(new_n370), .A3(new_n426), .A4(new_n429), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n295), .A2(new_n290), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n206), .A2(G33), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(G116), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G116), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n295), .A2(new_n434), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n289), .A2(new_n230), .B1(G20), .B2(new_n434), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G283), .ZN(new_n437));
  OAI211_X1 g0237(.A(new_n437), .B(new_n207), .C1(G33), .C2(new_n213), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n436), .A2(KEYINPUT20), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT20), .B1(new_n436), .B2(new_n438), .ZN(new_n440));
  OAI211_X1 g0240(.A(new_n433), .B(new_n435), .C1(new_n439), .C2(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(KEYINPUT83), .A2(G303), .ZN(new_n442));
  NAND2_X1  g0242(.A1(KEYINPUT83), .A2(G303), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n256), .A2(new_n442), .A3(new_n257), .A4(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(G264), .B(G1698), .C1(new_n251), .C2(new_n252), .ZN(new_n445));
  OAI211_X1 g0245(.A(G257), .B(new_n250), .C1(new_n251), .C2(new_n252), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n269), .ZN(new_n448));
  INV_X1    g0248(.A(G41), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n449), .A2(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(KEYINPUT5), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n450), .A2(new_n206), .A3(G45), .A4(new_n451), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n452), .A2(new_n272), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n452), .A2(G270), .A3(new_n268), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n448), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n441), .B1(new_n455), .B2(G200), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n448), .A2(new_n453), .A3(G190), .A4(new_n454), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT84), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n456), .A2(KEYINPUT84), .A3(new_n457), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n455), .A2(G169), .A3(new_n441), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT21), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n455), .A2(new_n338), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(new_n441), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n455), .A2(new_n441), .A3(KEYINPUT21), .A4(G169), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n465), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n258), .A2(new_n207), .A3(G87), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT85), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n472), .A2(KEYINPUT22), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT85), .B(KEYINPUT22), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n258), .A2(new_n475), .A3(new_n207), .A4(G87), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT23), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n207), .B2(G107), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n333), .A2(KEYINPUT23), .A3(G20), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n474), .A2(new_n476), .A3(new_n477), .A4(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT24), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n471), .A2(new_n473), .B1(new_n479), .B2(new_n480), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n485), .A2(KEYINPUT24), .A3(new_n476), .A4(new_n477), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n290), .A3(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n294), .A2(G107), .ZN(new_n488));
  OR2_X1    g0288(.A1(new_n488), .A2(KEYINPUT25), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT86), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n490), .B1(new_n488), .B2(KEYINPUT25), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n431), .A2(new_n432), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(new_n333), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n489), .A2(new_n491), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n487), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n258), .A2(G250), .A3(new_n250), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G294), .ZN(new_n499));
  OAI211_X1 g0299(.A(new_n498), .B(new_n499), .C1(new_n335), .C2(new_n214), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n269), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n452), .A2(new_n268), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(G264), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n501), .A2(new_n453), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(new_n338), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n500), .A2(new_n269), .B1(new_n502), .B2(G264), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(new_n453), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n346), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n497), .A2(new_n505), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n462), .A2(new_n470), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT82), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n206), .A2(G45), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n512), .B(G250), .C1(new_n267), .C2(new_n230), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n222), .A2(new_n250), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n212), .A2(G1698), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n515), .B(new_n516), .C1(new_n251), .C2(new_n252), .ZN(new_n517));
  NAND2_X1  g0317(.A1(G33), .A2(G116), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n514), .B1(new_n519), .B2(new_n269), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n512), .A2(new_n272), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT78), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n268), .B1(new_n517), .B2(new_n518), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT78), .ZN(new_n525));
  NOR4_X1   g0325(.A1(new_n524), .A2(new_n525), .A3(new_n514), .A4(new_n521), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n511), .B1(new_n527), .B2(new_n365), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n363), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n431), .A2(G87), .A3(new_n432), .ZN(new_n530));
  XNOR2_X1  g0330(.A(new_n530), .B(KEYINPUT81), .ZN(new_n531));
  INV_X1    g0331(.A(new_n324), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(new_n295), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT19), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n307), .B2(new_n213), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT79), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n258), .A2(new_n207), .A3(G68), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n207), .B1(new_n261), .B2(new_n534), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n372), .A2(new_n213), .A3(new_n333), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n537), .A2(new_n538), .A3(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n535), .A2(new_n536), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n290), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n531), .A2(new_n533), .A3(new_n544), .ZN(new_n545));
  OAI211_X1 g0345(.A(KEYINPUT82), .B(G190), .C1(new_n523), .C2(new_n526), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n528), .A2(new_n529), .A3(new_n545), .A4(new_n546), .ZN(new_n547));
  XNOR2_X1  g0347(.A(new_n324), .B(KEYINPUT80), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n544), .B(new_n533), .C1(new_n493), .C2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n338), .B1(new_n523), .B2(new_n526), .ZN(new_n551));
  INV_X1    g0351(.A(new_n527), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n550), .B(new_n551), .C1(new_n552), .C2(G169), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n547), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT77), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(KEYINPUT4), .ZN(new_n556));
  OAI211_X1 g0356(.A(G244), .B(new_n250), .C1(new_n251), .C2(new_n252), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n555), .A2(KEYINPUT4), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n334), .A2(G250), .ZN(new_n560));
  INV_X1    g0360(.A(new_n556), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n258), .A2(G244), .A3(new_n250), .A4(new_n561), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n559), .A2(new_n437), .A3(new_n560), .A4(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n269), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n502), .A2(G257), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n564), .A2(new_n453), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G200), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT6), .ZN(new_n568));
  NOR3_X1   g0368(.A1(new_n568), .A2(new_n213), .A3(G107), .ZN(new_n569));
  XNOR2_X1  g0369(.A(G97), .B(G107), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n569), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  OAI22_X1  g0371(.A1(new_n571), .A2(new_n207), .B1(new_n211), .B2(new_n352), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n397), .B1(new_n258), .B2(G20), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n262), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n333), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n290), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n295), .A2(new_n213), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n431), .A2(G97), .A3(new_n432), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n567), .B(new_n580), .C1(new_n365), .C2(new_n566), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n563), .A2(new_n269), .B1(G257), .B2(new_n502), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(new_n338), .A3(new_n453), .ZN(new_n583));
  INV_X1    g0383(.A(new_n566), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n583), .B(new_n579), .C1(new_n584), .C2(G169), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n507), .A2(G200), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n506), .A2(G190), .A3(new_n453), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n586), .A2(new_n487), .A3(new_n587), .A4(new_n496), .ZN(new_n588));
  NAND3_X1  g0388(.A1(new_n581), .A2(new_n585), .A3(new_n588), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n510), .A2(new_n554), .A3(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n430), .A2(new_n590), .ZN(G372));
  AND3_X1   g0391(.A1(new_n581), .A2(new_n585), .A3(new_n588), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n520), .A2(new_n522), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n363), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n545), .B(new_n594), .C1(new_n527), .C2(new_n365), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n346), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n551), .A2(new_n550), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n497), .A2(new_n508), .A3(new_n505), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n592), .B(new_n598), .C1(new_n599), .C2(new_n469), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT26), .ZN(new_n601));
  INV_X1    g0401(.A(new_n585), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n598), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(KEYINPUT26), .B1(new_n554), .B2(new_n585), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n600), .A2(new_n603), .A3(new_n597), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n430), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n318), .A2(new_n347), .A3(new_n344), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n425), .B1(new_n315), .B2(new_n607), .ZN(new_n608));
  AOI211_X1 g0408(.A(KEYINPUT87), .B(new_n386), .C1(new_n409), .C2(new_n410), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT87), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n610), .B1(new_n414), .B2(new_n415), .ZN(new_n611));
  NOR3_X1   g0411(.A1(new_n609), .A2(new_n611), .A3(new_n371), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n414), .A2(new_n415), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(KEYINPUT87), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n414), .A2(new_n610), .A3(new_n415), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT18), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n367), .B1(new_n608), .B2(new_n617), .ZN(new_n618));
  AND2_X1   g0418(.A1(new_n618), .A2(new_n369), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n606), .A2(new_n619), .ZN(G369));
  INV_X1    g0420(.A(G13), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n621), .A2(G20), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n206), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(G213), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(G343), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n497), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n599), .B1(new_n588), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n509), .A2(new_n628), .ZN(new_n631));
  INV_X1    g0431(.A(new_n628), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n469), .A2(new_n632), .ZN(new_n633));
  OR3_X1    g0433(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(new_n631), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n633), .B1(new_n630), .B2(new_n631), .ZN(new_n637));
  INV_X1    g0437(.A(G330), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n628), .A2(new_n441), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n462), .A2(new_n470), .A3(new_n639), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n469), .A2(new_n441), .A3(new_n628), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n637), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n636), .A2(new_n643), .ZN(G399));
  INV_X1    g0444(.A(new_n226), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n645), .A2(G41), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G1), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n540), .A2(G116), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n648), .A2(new_n649), .B1(new_n229), .B2(new_n647), .ZN(new_n650));
  XNOR2_X1  g0450(.A(new_n650), .B(KEYINPUT28), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n605), .A2(new_n632), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT29), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n598), .A2(new_n602), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT26), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n547), .A2(new_n553), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(new_n601), .A3(new_n602), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n597), .B(KEYINPUT91), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n655), .A2(new_n600), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(new_n632), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n660), .A2(KEYINPUT29), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n653), .A2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT88), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n566), .A2(new_n507), .A3(new_n663), .ZN(new_n664));
  OAI211_X1 g0464(.A(KEYINPUT88), .B(new_n453), .C1(new_n582), .C2(new_n506), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AND3_X1   g0466(.A1(new_n455), .A2(new_n593), .A3(new_n338), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n552), .A2(new_n582), .A3(new_n504), .A4(new_n466), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT30), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT89), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n669), .A2(new_n670), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n668), .A2(new_n671), .A3(KEYINPUT89), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  AND3_X1   g0477(.A1(new_n677), .A2(KEYINPUT31), .A3(new_n628), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n462), .A2(new_n470), .A3(new_n509), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n679), .A2(new_n656), .A3(new_n592), .A4(new_n632), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT90), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n668), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n666), .A2(KEYINPUT90), .A3(new_n667), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n682), .A2(new_n675), .A3(new_n671), .A4(new_n683), .ZN(new_n684));
  AOI22_X1  g0484(.A1(new_n680), .A2(KEYINPUT31), .B1(new_n684), .B2(new_n628), .ZN(new_n685));
  OAI21_X1  g0485(.A(G330), .B1(new_n678), .B2(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n662), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n651), .B1(new_n688), .B2(G1), .ZN(G364));
  INV_X1    g0489(.A(new_n642), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n648), .B1(G45), .B2(new_n622), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n640), .A2(new_n638), .A3(new_n641), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT92), .Z(new_n695));
  NOR3_X1   g0495(.A1(G13), .A2(G20), .A3(G33), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n640), .A2(new_n641), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n645), .A2(new_n258), .ZN(new_n698));
  INV_X1    g0498(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n699), .B1(new_n244), .B2(G45), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(G45), .B2(new_n229), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n226), .A2(G355), .A3(new_n258), .ZN(new_n702));
  OAI211_X1 g0502(.A(new_n701), .B(new_n702), .C1(G116), .C2(new_n226), .ZN(new_n703));
  AND2_X1   g0503(.A1(KEYINPUT93), .A2(G169), .ZN(new_n704));
  NOR2_X1   g0504(.A1(KEYINPUT93), .A2(G169), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n230), .B1(new_n706), .B2(G20), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(new_n696), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n207), .A2(new_n365), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n338), .A2(new_n418), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n338), .A2(G200), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI22_X1  g0516(.A1(G326), .A2(new_n713), .B1(new_n716), .B2(G322), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n207), .A2(G190), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n711), .A2(new_n718), .ZN(new_n719));
  XOR2_X1   g0519(.A(KEYINPUT33), .B(G317), .Z(new_n720));
  OAI211_X1 g0520(.A(new_n717), .B(new_n262), .C1(new_n719), .C2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n363), .A2(new_n338), .A3(new_n710), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n721), .B1(G303), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G179), .A2(G200), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G190), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(G294), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n718), .A2(new_n714), .A3(KEYINPUT94), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT94), .B1(new_n718), .B2(new_n714), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G311), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n718), .A2(new_n725), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n734), .A2(KEYINPUT97), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(KEYINPUT97), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n363), .A2(new_n338), .A3(new_n718), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n738), .A2(G329), .B1(G283), .B2(new_n740), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n724), .A2(new_n728), .A3(new_n733), .A4(new_n741), .ZN(new_n742));
  OR2_X1    g0542(.A1(new_n731), .A2(KEYINPUT95), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n731), .A2(KEYINPUT95), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G77), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n740), .A2(G107), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n734), .A2(new_n393), .ZN(new_n749));
  XOR2_X1   g0549(.A(KEYINPUT96), .B(KEYINPUT32), .Z(new_n750));
  XOR2_X1   g0550(.A(new_n749), .B(new_n750), .Z(new_n751));
  INV_X1    g0551(.A(new_n719), .ZN(new_n752));
  AOI22_X1  g0552(.A1(new_n752), .A2(G68), .B1(new_n727), .B2(G97), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(new_n400), .B2(new_n715), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n722), .A2(new_n372), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n754), .A2(new_n262), .A3(new_n755), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n747), .A2(new_n748), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n712), .A2(new_n202), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n742), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n707), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n697), .A2(new_n709), .A3(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n695), .B1(new_n692), .B2(new_n761), .ZN(G396));
  OAI21_X1  g0562(.A(new_n428), .B1(new_n330), .B2(new_n632), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n348), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n344), .A2(new_n347), .A3(new_n632), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n652), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n766), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n768), .A2(new_n605), .A3(new_n632), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n687), .B(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n692), .ZN(new_n772));
  NOR2_X1   g0572(.A1(G13), .A2(G33), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n766), .A2(new_n773), .ZN(new_n774));
  AOI22_X1  g0574(.A1(G143), .A2(new_n716), .B1(new_n752), .B2(G150), .ZN(new_n775));
  INV_X1    g0575(.A(G137), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n775), .B1(new_n776), .B2(new_n712), .C1(new_n745), .C2(new_n393), .ZN(new_n777));
  XNOR2_X1  g0577(.A(new_n777), .B(KEYINPUT34), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n739), .A2(new_n221), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n258), .B1(new_n722), .B2(new_n202), .ZN(new_n780));
  AOI211_X1 g0580(.A(new_n779), .B(new_n780), .C1(G58), .C2(new_n727), .ZN(new_n781));
  INV_X1    g0581(.A(G132), .ZN(new_n782));
  OAI211_X1 g0582(.A(new_n778), .B(new_n781), .C1(new_n782), .C2(new_n737), .ZN(new_n783));
  INV_X1    g0583(.A(G311), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n737), .A2(new_n784), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n746), .A2(G116), .B1(G97), .B2(new_n727), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n740), .A2(G87), .B1(G283), .B2(new_n752), .ZN(new_n787));
  INV_X1    g0587(.A(G294), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n262), .B1(new_n715), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n722), .A2(new_n333), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n789), .B(new_n790), .C1(G303), .C2(new_n713), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n786), .A2(new_n787), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n783), .B1(new_n785), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(new_n707), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n707), .A2(new_n773), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(new_n211), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n774), .A2(new_n691), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n772), .A2(new_n797), .ZN(G384));
  AND3_X1   g0598(.A1(new_n684), .A2(KEYINPUT31), .A3(new_n628), .ZN(new_n799));
  OAI21_X1  g0599(.A(KEYINPUT103), .B1(new_n685), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(KEYINPUT103), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n684), .A2(KEYINPUT31), .A3(new_n628), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT31), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(new_n590), .B2(new_n632), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n684), .A2(new_n628), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n801), .B(new_n802), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n800), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n319), .A2(new_n321), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n314), .B(new_n628), .C1(new_n808), .C2(new_n288), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n315), .B(new_n318), .C1(new_n313), .C2(new_n632), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n807), .A2(new_n768), .A3(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT38), .ZN(new_n813));
  INV_X1    g0613(.A(new_n626), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n414), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT37), .ZN(new_n816));
  NAND4_X1  g0616(.A1(new_n613), .A2(new_n815), .A3(new_n816), .A4(new_n421), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n609), .A2(new_n611), .ZN(new_n819));
  INV_X1    g0619(.A(new_n421), .ZN(new_n820));
  OAI21_X1  g0620(.A(KEYINPUT99), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT99), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n822), .B(new_n421), .C1(new_n609), .C2(new_n611), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n821), .A2(new_n815), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n818), .B1(new_n824), .B2(KEYINPUT37), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT100), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n425), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n423), .A2(KEYINPUT100), .A3(new_n424), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n827), .B(new_n828), .C1(new_n612), .C2(new_n616), .ZN(new_n829));
  INV_X1    g0629(.A(new_n815), .ZN(new_n830));
  AND2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n813), .B1(new_n825), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n407), .A2(new_n389), .ZN(new_n833));
  OAI211_X1 g0633(.A(new_n814), .B(new_n833), .C1(new_n417), .C2(new_n425), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n386), .A2(new_n626), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n820), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n817), .B1(new_n836), .B2(new_n816), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n834), .A2(new_n837), .A3(KEYINPUT38), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n812), .B1(new_n832), .B2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT98), .ZN(new_n840));
  AND3_X1   g0640(.A1(new_n834), .A2(new_n837), .A3(KEYINPUT38), .ZN(new_n841));
  AOI21_X1  g0641(.A(KEYINPUT38), .B1(new_n834), .B2(new_n837), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n840), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n834), .A2(new_n837), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n813), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(KEYINPUT98), .A3(new_n838), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n766), .B1(new_n800), .B2(new_n806), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n843), .A2(new_n846), .A3(new_n847), .A4(new_n811), .ZN(new_n848));
  XOR2_X1   g0648(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n849));
  AOI22_X1  g0649(.A1(new_n839), .A2(KEYINPUT40), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AND2_X1   g0650(.A1(new_n430), .A2(new_n807), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n823), .A2(new_n815), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n614), .A2(new_n615), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n822), .B1(new_n854), .B2(new_n421), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT37), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  AOI22_X1  g0656(.A1(new_n856), .A2(new_n817), .B1(new_n830), .B2(new_n829), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n838), .B1(new_n857), .B2(KEYINPUT38), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n807), .A2(new_n768), .A3(new_n811), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(new_n859), .A3(KEYINPUT40), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n843), .A2(new_n846), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n849), .B1(new_n861), .B2(new_n812), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n862), .A3(G330), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n430), .A2(G330), .A3(new_n807), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n852), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n866), .B(KEYINPUT101), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n662), .A2(new_n430), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n619), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n867), .B(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n617), .A2(new_n626), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n769), .A2(new_n765), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n811), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n871), .B1(new_n861), .B2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT39), .ZN(new_n875));
  NOR3_X1   g0675(.A1(new_n841), .A2(new_n842), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n876), .B1(new_n858), .B2(new_n875), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n288), .A2(new_n314), .A3(new_n632), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n874), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n870), .B(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n881), .B1(new_n206), .B2(new_n622), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT35), .ZN(new_n883));
  AOI211_X1 g0683(.A(new_n207), .B(new_n230), .C1(new_n571), .C2(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(new_n884), .B(G116), .C1(new_n883), .C2(new_n571), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT36), .ZN(new_n886));
  OAI21_X1  g0686(.A(G77), .B1(new_n400), .B2(new_n221), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n887), .A2(new_n229), .B1(G50), .B2(new_n221), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n888), .A2(G1), .A3(new_n621), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n882), .A2(new_n886), .A3(new_n889), .ZN(G367));
  OAI211_X1 g0690(.A(new_n581), .B(new_n585), .C1(new_n580), .C2(new_n632), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n602), .A2(new_n628), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n634), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT42), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n585), .B1(new_n891), .B2(new_n509), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n897), .A2(new_n632), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n598), .B1(new_n545), .B2(new_n632), .ZN(new_n900));
  OR3_X1    g0700(.A1(new_n597), .A2(new_n545), .A3(new_n632), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OR3_X1    g0702(.A1(new_n899), .A2(KEYINPUT43), .A3(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n643), .A2(new_n894), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n902), .A2(KEYINPUT43), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n902), .A2(KEYINPUT43), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n899), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n903), .A2(new_n904), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n903), .A2(new_n908), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n910), .B1(new_n643), .B2(new_n894), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n646), .B(KEYINPUT41), .ZN(new_n912));
  INV_X1    g0712(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n642), .B1(new_n634), .B2(new_n637), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT105), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT105), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n643), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n915), .B1(new_n914), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT44), .B1(new_n636), .B2(new_n893), .ZN(new_n919));
  XOR2_X1   g0719(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n920));
  NAND3_X1  g0720(.A1(new_n636), .A2(new_n893), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n634), .A2(new_n635), .ZN(new_n922));
  INV_X1    g0722(.A(KEYINPUT44), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n922), .A2(new_n923), .A3(new_n894), .ZN(new_n924));
  INV_X1    g0724(.A(new_n920), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n922), .B2(new_n894), .ZN(new_n926));
  NAND4_X1  g0726(.A1(new_n919), .A2(new_n921), .A3(new_n924), .A4(new_n926), .ZN(new_n927));
  NAND4_X1  g0727(.A1(new_n688), .A2(KEYINPUT106), .A3(new_n918), .A4(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT106), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n918), .A2(new_n686), .A3(new_n661), .A4(new_n653), .ZN(new_n930));
  AND4_X1   g0730(.A1(new_n919), .A2(new_n921), .A3(new_n924), .A4(new_n926), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n913), .B1(new_n933), .B2(new_n688), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n206), .B1(new_n622), .B2(G45), .ZN(new_n935));
  INV_X1    g0735(.A(new_n935), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n909), .B(new_n911), .C1(new_n934), .C2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n727), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n938), .A2(new_n221), .ZN(new_n939));
  INV_X1    g0739(.A(new_n939), .ZN(new_n940));
  AOI22_X1  g0740(.A1(G143), .A2(new_n713), .B1(new_n716), .B2(G150), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT107), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n745), .A2(new_n202), .B1(new_n393), .B2(new_n719), .ZN(new_n943));
  XOR2_X1   g0743(.A(new_n943), .B(KEYINPUT108), .Z(new_n944));
  NAND3_X1  g0744(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT107), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n945), .B1(new_n400), .B2(new_n722), .C1(new_n211), .C2(new_n739), .ZN(new_n946));
  OR3_X1    g0746(.A1(new_n944), .A2(new_n262), .A3(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n734), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n942), .B(new_n947), .C1(G137), .C2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n746), .A2(G283), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n948), .A2(G317), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n740), .A2(G97), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n950), .A2(new_n262), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n938), .A2(new_n333), .B1(new_n719), .B2(new_n788), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n442), .A2(new_n443), .ZN(new_n955));
  OAI22_X1  g0755(.A1(new_n712), .A2(new_n784), .B1(new_n715), .B2(new_n955), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n953), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n723), .A2(G116), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT46), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n949), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(KEYINPUT47), .Z(new_n961));
  NAND2_X1  g0761(.A1(new_n961), .A2(new_n707), .ZN(new_n962));
  OAI221_X1 g0762(.A(new_n708), .B1(new_n226), .B2(new_n532), .C1(new_n699), .C2(new_n240), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n900), .A2(new_n696), .A3(new_n901), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n962), .A2(new_n691), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n937), .A2(new_n965), .ZN(G387));
  INV_X1    g0766(.A(new_n918), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n662), .B2(new_n687), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n968), .A2(new_n646), .A3(new_n930), .ZN(new_n969));
  INV_X1    g0769(.A(G317), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n784), .A2(new_n719), .B1(new_n715), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G322), .B2(new_n713), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n972), .B1(new_n745), .B2(new_n955), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(KEYINPUT48), .ZN(new_n974));
  INV_X1    g0774(.A(G283), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n974), .B1(new_n975), .B2(new_n938), .C1(new_n788), .C2(new_n722), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT49), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n740), .A2(G116), .B1(G326), .B2(new_n948), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n977), .A2(new_n262), .A3(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n732), .A2(G68), .B1(G97), .B2(new_n740), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n351), .B2(new_n734), .C1(new_n387), .C2(new_n719), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G50), .B2(new_n716), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n548), .A2(new_n727), .ZN(new_n983));
  OAI211_X1 g0783(.A(new_n982), .B(new_n983), .C1(new_n393), .C2(new_n712), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n723), .A2(G77), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n258), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n979), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n707), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n696), .B1(new_n630), .B2(new_n631), .ZN(new_n989));
  INV_X1    g0789(.A(G45), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n698), .B1(new_n236), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n226), .A2(new_n649), .A3(new_n258), .ZN(new_n992));
  AOI211_X1 g0792(.A(G45), .B(new_n649), .C1(G68), .C2(G77), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n387), .A2(G50), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT50), .ZN(new_n995));
  AOI22_X1  g0795(.A1(new_n991), .A2(new_n992), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n226), .A2(G107), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n708), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n988), .A2(new_n989), .A3(new_n998), .ZN(new_n999));
  OAI221_X1 g0799(.A(new_n969), .B1(new_n935), .B2(new_n967), .C1(new_n692), .C2(new_n999), .ZN(G393));
  INV_X1    g0800(.A(KEYINPUT112), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n643), .A2(KEYINPUT109), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n643), .A2(KEYINPUT109), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n931), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n927), .A2(KEYINPUT109), .A3(new_n643), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n935), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n894), .A2(new_n696), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n258), .B1(new_n948), .B2(G322), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n748), .B(new_n1009), .C1(new_n434), .C2(new_n938), .ZN(new_n1010));
  OAI22_X1  g0810(.A1(new_n712), .A2(new_n970), .B1(new_n715), .B2(new_n784), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT52), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n1010), .A2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n723), .A2(G283), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n732), .A2(G294), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n719), .A2(new_n955), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n740), .A2(G87), .B1(G143), .B2(new_n948), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n1020), .B(new_n258), .C1(new_n221), .C2(new_n722), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT111), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n727), .A2(G77), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n746), .A2(new_n327), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n712), .A2(new_n351), .B1(new_n715), .B2(new_n393), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT51), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1025), .A2(new_n1026), .B1(G50), .B2(new_n752), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1022), .A2(new_n1023), .A3(new_n1024), .A4(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1019), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n707), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n708), .B1(new_n213), .B2(new_n226), .C1(new_n699), .C2(new_n248), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n691), .A2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT110), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1008), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1001), .B1(new_n1007), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1006), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1002), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n927), .A2(new_n1039), .A3(new_n1003), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  OAI211_X1 g0841(.A(KEYINPUT112), .B(new_n1035), .C1(new_n1041), .C2(new_n935), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n1041), .A2(new_n930), .B1(new_n932), .B2(new_n928), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n1037), .A2(new_n1042), .B1(new_n1043), .B2(new_n646), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(G390));
  NAND2_X1  g0845(.A1(new_n873), .A2(new_n878), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n877), .A2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n829), .A2(new_n830), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n823), .A2(new_n815), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n816), .B1(new_n1050), .B2(new_n821), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1049), .B1(new_n1051), .B2(new_n818), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n841), .B1(new_n1052), .B2(new_n813), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n659), .A2(new_n632), .A3(new_n764), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n765), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n809), .A2(new_n810), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n878), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1053), .A2(new_n1058), .ZN(new_n1059));
  OAI211_X1 g0859(.A(G330), .B(new_n859), .C1(new_n1048), .C2(new_n1059), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n687), .A2(new_n768), .A3(new_n811), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n1061), .B1(new_n1053), .B2(new_n1058), .C1(new_n877), .C2(new_n1047), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n936), .A3(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n877), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n773), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n692), .B1(new_n795), .B2(new_n387), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n258), .B1(new_n715), .B2(new_n782), .ZN(new_n1068));
  XOR2_X1   g0868(.A(KEYINPUT54), .B(G143), .Z(new_n1069));
  AOI21_X1  g0869(.A(new_n1068), .B1(new_n746), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(G128), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1070), .B1(new_n1071), .B2(new_n712), .C1(new_n776), .C2(new_n719), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n739), .A2(new_n202), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n723), .A2(G150), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT53), .ZN(new_n1075));
  INV_X1    g0875(.A(G125), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n737), .A2(new_n1076), .B1(new_n393), .B2(new_n938), .ZN(new_n1077));
  NOR4_X1   g0877(.A1(new_n1072), .A2(new_n1073), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1023), .B1(new_n975), .B2(new_n712), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n755), .B(new_n1079), .C1(new_n738), .C2(G294), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n262), .B1(new_n715), .B2(new_n434), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n1081), .B(new_n779), .C1(G107), .C2(new_n752), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1083), .B1(G97), .B2(new_n746), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n707), .B1(new_n1078), .B2(new_n1084), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1066), .A2(KEYINPUT113), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1065), .A2(new_n1067), .A3(new_n1085), .A4(new_n1086), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n868), .A2(new_n864), .A3(new_n619), .ZN(new_n1088));
  AND2_X1   g0888(.A1(new_n847), .A2(G330), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1061), .B(new_n1056), .C1(new_n1089), .C2(new_n811), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1057), .B1(new_n686), .B2(new_n766), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n812), .B2(new_n638), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n872), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1088), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n1059), .B1(new_n1064), .B2(new_n1046), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n859), .A2(G330), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1062), .B(new_n1094), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(new_n646), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1094), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1063), .B(new_n1087), .C1(new_n1098), .C2(new_n1099), .ZN(G378));
  NAND2_X1  g0900(.A1(new_n355), .A2(new_n814), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n370), .B(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1103));
  XOR2_X1   g0903(.A(new_n1102), .B(new_n1103), .Z(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n863), .B2(KEYINPUT118), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT118), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n860), .A2(new_n862), .A3(new_n1106), .A4(G330), .ZN(new_n1107));
  AND2_X1   g0907(.A1(new_n880), .A2(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n880), .A2(new_n1107), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1105), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n863), .A2(KEYINPUT118), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1104), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n876), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n879), .B(new_n1114), .C1(new_n1053), .C2(KEYINPUT39), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n843), .A2(new_n846), .A3(new_n872), .A4(new_n811), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n1116), .A2(new_n871), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n1118), .A2(new_n850), .A3(new_n1106), .A4(G330), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n880), .A2(new_n1107), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1113), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1110), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1088), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1123), .A2(KEYINPUT120), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(KEYINPUT120), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1097), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1122), .A2(KEYINPUT57), .A3(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(KEYINPUT121), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT57), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT121), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1122), .A2(new_n1132), .A3(new_n1126), .A4(KEYINPUT57), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1128), .A2(new_n1131), .A3(new_n646), .A4(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n712), .A2(new_n434), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1135), .B(new_n939), .C1(G107), .C2(new_n716), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n740), .A2(G58), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1136), .A2(new_n449), .A3(new_n1137), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n732), .A2(new_n548), .B1(G97), .B2(new_n752), .ZN(new_n1139));
  OR2_X1    g0939(.A1(new_n1139), .A2(KEYINPUT114), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(KEYINPUT114), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1140), .A2(new_n262), .A3(new_n985), .A4(new_n1141), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1138), .B(new_n1142), .C1(G283), .C2(new_n738), .ZN(new_n1143));
  XNOR2_X1  g0943(.A(new_n1143), .B(KEYINPUT115), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT58), .Z(new_n1145));
  OAI21_X1  g0945(.A(new_n202), .B1(new_n251), .B2(G41), .ZN(new_n1146));
  AOI21_X1  g0946(.A(G33), .B1(new_n948), .B2(G124), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1147), .B(new_n449), .C1(new_n393), .C2(new_n739), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT117), .ZN(new_n1149));
  OAI22_X1  g0949(.A1(new_n731), .A2(new_n776), .B1(new_n1076), .B2(new_n712), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n723), .A2(new_n1069), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT116), .ZN(new_n1152));
  AOI211_X1 g0952(.A(new_n1150), .B(new_n1152), .C1(G128), .C2(new_n716), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n1153), .B1(new_n782), .B2(new_n719), .C1(new_n351), .C2(new_n938), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT59), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1145), .B(new_n1146), .C1(new_n1149), .C2(new_n1155), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1156), .A2(new_n707), .B1(new_n202), .B2(new_n795), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n691), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1158), .B1(new_n773), .B2(new_n1104), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(new_n1122), .B2(new_n936), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT119), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n935), .B1(new_n1110), .B2(new_n1121), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT119), .B1(new_n1163), .B2(new_n1159), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1162), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1134), .A2(new_n1165), .ZN(G375));
  INV_X1    g0966(.A(new_n1094), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1090), .A2(new_n1093), .A3(new_n1088), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1167), .A2(new_n912), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n935), .B1(new_n1090), .B2(new_n1093), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1057), .A2(new_n773), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n738), .A2(G303), .B1(G294), .B2(new_n713), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1172), .B1(new_n211), .B2(new_n739), .C1(new_n434), .C2(new_n719), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n745), .A2(new_n333), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n715), .A2(new_n975), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n983), .B(new_n262), .C1(new_n213), .C2(new_n722), .ZN(new_n1176));
  NOR4_X1   g0976(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n723), .A2(G159), .B1(G50), .B2(new_n727), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n713), .A2(G132), .B1(new_n752), .B2(new_n1069), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1178), .A2(new_n258), .A3(new_n1179), .ZN(new_n1180));
  OAI221_X1 g0980(.A(new_n1137), .B1(new_n731), .B2(new_n351), .C1(new_n1071), .C2(new_n737), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1180), .B(new_n1181), .C1(G137), .C2(new_n716), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n707), .B1(new_n1177), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n795), .A2(new_n221), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1171), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1170), .B1(new_n691), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1169), .A2(new_n1186), .ZN(G381));
  INV_X1    g0987(.A(G378), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1134), .A2(new_n1188), .A3(new_n1165), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1189), .A2(G384), .A3(G381), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1044), .A2(new_n937), .A3(new_n965), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1191), .A2(G396), .A3(G393), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1190), .A2(new_n1192), .ZN(G407));
  OAI211_X1 g0993(.A(G407), .B(G213), .C1(G343), .C2(new_n1189), .ZN(G409));
  INV_X1    g0994(.A(KEYINPUT122), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT60), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1168), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1197), .A2(new_n646), .A3(new_n1167), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1196), .B1(new_n1168), .B2(new_n1195), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1186), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n772), .A3(new_n797), .ZN(new_n1201));
  OAI211_X1 g1001(.A(G384), .B(new_n1186), .C1(new_n1198), .C2(new_n1199), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n627), .A2(G213), .ZN(new_n1203));
  OR2_X1    g1003(.A1(new_n1203), .A2(KEYINPUT123), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1201), .A2(new_n1202), .A3(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n627), .A2(G213), .A3(G2897), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  XNOR2_X1  g1007(.A(new_n1205), .B(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(G375), .A2(G378), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1122), .A2(new_n912), .A3(new_n1126), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1188), .A2(new_n1160), .A3(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1211), .A2(new_n1203), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1208), .B1(new_n1209), .B2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1188), .B1(new_n1134), .B2(new_n1165), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1216));
  NOR3_X1   g1016(.A1(new_n1215), .A2(new_n1212), .A3(new_n1216), .ZN(new_n1217));
  OAI21_X1  g1017(.A(KEYINPUT63), .B1(new_n1214), .B2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1212), .B1(G375), .B2(G378), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1216), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT63), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  XOR2_X1   g1023(.A(G393), .B(G396), .Z(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1191), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1044), .B1(new_n937), .B2(new_n965), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1225), .B1(new_n1226), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT125), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  OAI211_X1 g1030(.A(KEYINPUT125), .B(new_n1225), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1230), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(G387), .A2(G390), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n1233), .A2(new_n1191), .A3(new_n1224), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(KEYINPUT124), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT124), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1233), .A2(new_n1236), .A3(new_n1191), .A4(new_n1224), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1235), .A2(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1232), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT61), .ZN(new_n1240));
  AOI21_X1  g1040(.A(KEYINPUT126), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT126), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1242), .B(KEYINPUT61), .C1(new_n1232), .C2(new_n1238), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1241), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1218), .A2(new_n1223), .A3(new_n1244), .ZN(new_n1245));
  XOR2_X1   g1045(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1246));
  OAI21_X1  g1046(.A(new_n1246), .B1(new_n1219), .B2(new_n1208), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT62), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(new_n1215), .A2(new_n1212), .A3(KEYINPUT62), .A4(new_n1216), .ZN(new_n1250));
  NOR3_X1   g1050(.A1(new_n1247), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1245), .B1(new_n1251), .B2(new_n1239), .ZN(G405));
  INV_X1    g1052(.A(new_n1189), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1220), .B1(new_n1253), .B2(new_n1215), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1209), .A2(new_n1189), .A3(new_n1216), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(new_n1239), .ZN(G402));
endmodule


