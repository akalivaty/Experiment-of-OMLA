//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 0 0 1 1 1 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 1 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034;
  INV_X1    g000(.A(G116), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT67), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G116), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n188), .A2(new_n190), .A3(G119), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G116), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT68), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT69), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT2), .B(G113), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n191), .A2(KEYINPUT68), .A3(new_n193), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n196), .A2(new_n197), .A3(new_n198), .A4(new_n199), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n191), .A2(KEYINPUT68), .A3(new_n193), .ZN(new_n201));
  AOI21_X1  g015(.A(KEYINPUT68), .B1(new_n191), .B2(new_n193), .ZN(new_n202));
  INV_X1    g016(.A(new_n198), .ZN(new_n203));
  NOR3_X1   g017(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n203), .A2(new_n191), .A3(new_n193), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT69), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n200), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  INV_X1    g024(.A(G128), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n212));
  INV_X1    g026(.A(G146), .ZN(new_n213));
  AND3_X1   g027(.A1(new_n213), .A2(KEYINPUT65), .A3(G143), .ZN(new_n214));
  AOI21_X1  g028(.A(KEYINPUT65), .B1(new_n213), .B2(G143), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n210), .B(new_n212), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  NOR2_X1   g030(.A1(new_n209), .A2(G146), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT64), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n218), .B1(new_n213), .B2(G143), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n209), .A2(KEYINPUT64), .A3(G146), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n217), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n213), .A2(G143), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n211), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n216), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT11), .ZN(new_n225));
  INV_X1    g039(.A(G134), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n225), .B1(new_n226), .B2(G137), .ZN(new_n227));
  INV_X1    g041(.A(G137), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(KEYINPUT11), .A3(G134), .ZN(new_n229));
  INV_X1    g043(.A(G131), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n226), .A2(G137), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n227), .A2(new_n229), .A3(new_n230), .A4(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT66), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n226), .B2(G137), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n228), .A2(KEYINPUT66), .A3(G134), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n234), .A2(new_n231), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G131), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n224), .A2(new_n232), .A3(new_n237), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n209), .A2(KEYINPUT64), .A3(G146), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT64), .B1(new_n209), .B2(G146), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n222), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AND2_X1   g055(.A1(KEYINPUT0), .A2(G128), .ZN(new_n242));
  NOR2_X1   g056(.A1(KEYINPUT0), .A2(G128), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n213), .A2(G143), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT65), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n209), .B2(G146), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n213), .A2(KEYINPUT65), .A3(G143), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI22_X1  g063(.A1(new_n241), .A2(new_n244), .B1(new_n249), .B2(new_n242), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n227), .A2(new_n229), .A3(new_n231), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G131), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n232), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n238), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n255), .B1(new_n238), .B2(new_n254), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n208), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n237), .A2(new_n232), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n260), .A2(new_n224), .B1(new_n250), .B2(new_n253), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n207), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n263));
  INV_X1    g077(.A(G210), .ZN(new_n264));
  NOR3_X1   g078(.A1(new_n264), .A2(G237), .A3(G953), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n263), .B(new_n265), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT26), .B(G101), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n258), .A2(new_n262), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT31), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n258), .A2(KEYINPUT31), .A3(new_n262), .A4(new_n268), .ZN(new_n272));
  AND2_X1   g086(.A1(new_n252), .A2(new_n232), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n210), .B(new_n242), .C1(new_n214), .C2(new_n215), .ZN(new_n274));
  INV_X1    g088(.A(new_n244), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n274), .B1(new_n221), .B2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n223), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n241), .A2(new_n277), .B1(new_n249), .B2(new_n212), .ZN(new_n278));
  OAI22_X1  g092(.A1(new_n273), .A2(new_n276), .B1(new_n278), .B2(new_n259), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n280), .A2(KEYINPUT69), .A3(new_n205), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n279), .B1(new_n281), .B2(new_n200), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n207), .A2(new_n261), .ZN(new_n283));
  OAI21_X1  g097(.A(KEYINPUT28), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT28), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n262), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n268), .B(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(new_n289), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n271), .A2(new_n272), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(G472), .A2(G902), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT32), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n286), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n279), .A2(new_n281), .A3(new_n200), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n285), .B1(new_n262), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n290), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n279), .A2(KEYINPUT30), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n238), .A2(new_n254), .A3(new_n255), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n282), .B1(new_n301), .B2(new_n208), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT31), .B1(new_n302), .B2(new_n268), .ZN(new_n303));
  INV_X1    g117(.A(new_n272), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n298), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT32), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n306), .A3(new_n292), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n262), .B2(new_n285), .ZN(new_n309));
  AOI211_X1 g123(.A(KEYINPUT73), .B(KEYINPUT28), .C1(new_n207), .C2(new_n261), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n268), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT29), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT72), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n297), .A2(new_n315), .ZN(new_n316));
  AOI211_X1 g130(.A(KEYINPUT72), .B(new_n285), .C1(new_n262), .C2(new_n296), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n311), .B(new_n314), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n284), .A2(new_n286), .A3(new_n289), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n207), .B1(new_n299), .B2(new_n300), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n312), .B1(new_n320), .B2(new_n282), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n313), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G902), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n318), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n294), .A2(new_n307), .B1(G472), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(G952), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(G953), .ZN(new_n327));
  NAND2_X1  g141(.A1(G234), .A2(G237), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(G902), .A3(G953), .ZN(new_n331));
  INV_X1    g145(.A(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT21), .B(G898), .ZN(new_n333));
  AOI21_X1  g147(.A(new_n330), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(G214), .B1(G237), .B2(G902), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT87), .ZN(new_n338));
  OAI21_X1  g152(.A(G113), .B1(new_n193), .B2(KEYINPUT5), .ZN(new_n339));
  INV_X1    g153(.A(new_n193), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT67), .B(G116), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n340), .B1(new_n341), .B2(G119), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n339), .B1(new_n342), .B2(KEYINPUT5), .ZN(new_n343));
  INV_X1    g157(.A(new_n205), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n338), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT5), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n194), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g161(.A(KEYINPUT87), .B(new_n205), .C1(new_n347), .C2(new_n339), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(KEYINPUT82), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(KEYINPUT82), .ZN(new_n351));
  INV_X1    g165(.A(G107), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G104), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n350), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G101), .ZN(new_n355));
  INV_X1    g169(.A(G104), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(G107), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n349), .A2(new_n352), .A3(KEYINPUT82), .A4(G104), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n354), .A2(new_n355), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT83), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n360), .B1(new_n352), .B2(G104), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n353), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n357), .A2(new_n360), .ZN(new_n363));
  OAI21_X1  g177(.A(G101), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n359), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n345), .A2(new_n348), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n359), .A2(new_n364), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n346), .B1(new_n196), .B2(new_n199), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n367), .B(new_n205), .C1(new_n368), .C2(new_n339), .ZN(new_n369));
  XNOR2_X1  g183(.A(G110), .B(G122), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT8), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n366), .A2(new_n369), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(KEYINPUT88), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT88), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n366), .A2(new_n369), .A3(new_n374), .A4(new_n371), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n365), .B(new_n205), .C1(new_n368), .C2(new_n339), .ZN(new_n377));
  INV_X1    g191(.A(new_n354), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n358), .A2(new_n357), .ZN(new_n379));
  OAI21_X1  g193(.A(G101), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(KEYINPUT4), .A3(new_n359), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT4), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n382), .B(G101), .C1(new_n378), .C2(new_n379), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n377), .B(new_n370), .C1(new_n207), .C2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G125), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n278), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n276), .A2(G125), .ZN(new_n388));
  INV_X1    g202(.A(G224), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(G953), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT7), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AND3_X1   g206(.A1(new_n387), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n392), .B1(new_n387), .B2(new_n388), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  AND2_X1   g209(.A1(new_n385), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(G902), .B1(new_n376), .B2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n377), .B1(new_n207), .B2(new_n384), .ZN(new_n398));
  INV_X1    g212(.A(new_n370), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT6), .A3(new_n385), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT6), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n398), .A2(new_n402), .A3(new_n399), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n387), .A2(new_n388), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n404), .B(new_n390), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n401), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(G210), .B1(G237), .B2(G902), .ZN(new_n407));
  AND3_X1   g221(.A1(new_n397), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(new_n407), .B1(new_n397), .B2(new_n406), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n337), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT74), .B(G217), .ZN(new_n411));
  INV_X1    g225(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(G234), .B2(new_n323), .ZN(new_n413));
  XOR2_X1   g227(.A(new_n413), .B(KEYINPUT75), .Z(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT76), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(KEYINPUT79), .A2(KEYINPUT25), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT23), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n419), .B1(new_n192), .B2(G128), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n211), .A2(KEYINPUT23), .A3(G119), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n420), .B(new_n421), .C1(G119), .C2(new_n211), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G110), .ZN(new_n423));
  XOR2_X1   g237(.A(KEYINPUT24), .B(G110), .Z(new_n424));
  XNOR2_X1  g238(.A(G119), .B(G128), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n423), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(G140), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G125), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n386), .A2(G140), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT77), .A4(KEYINPUT16), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n429), .A2(new_n430), .A3(KEYINPUT16), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT16), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n428), .A3(G125), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT77), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n213), .B(new_n431), .C1(new_n432), .C2(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n429), .A2(new_n430), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n435), .B(new_n434), .C1(new_n439), .C2(new_n433), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n213), .B1(new_n440), .B2(new_n431), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n427), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n431), .B1(new_n432), .B2(new_n436), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(G146), .ZN(new_n444));
  OAI22_X1  g258(.A1(new_n422), .A2(G110), .B1(new_n425), .B2(new_n424), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n429), .A2(new_n430), .A3(new_n213), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G953), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(G221), .A3(G234), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n450), .B(KEYINPUT78), .ZN(new_n451));
  XNOR2_X1  g265(.A(KEYINPUT22), .B(G137), .ZN(new_n452));
  XOR2_X1   g266(.A(new_n451), .B(new_n452), .Z(new_n453));
  NAND2_X1  g267(.A1(new_n448), .A2(new_n453), .ZN(new_n454));
  XNOR2_X1  g268(.A(new_n451), .B(new_n452), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n442), .A2(new_n447), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n418), .B1(new_n457), .B2(new_n323), .ZN(new_n458));
  AOI211_X1 g272(.A(G902), .B(new_n417), .C1(new_n454), .C2(new_n456), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n416), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n457), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n414), .A2(new_n323), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n460), .A2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(G237), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n449), .A3(G214), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(KEYINPUT89), .B2(new_n209), .ZN(new_n468));
  XNOR2_X1  g282(.A(KEYINPUT89), .B(G143), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n468), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n470), .A2(G131), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT17), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n468), .B(new_n230), .C1(new_n467), .C2(new_n469), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(KEYINPUT17), .A3(G131), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n474), .A2(new_n437), .A3(new_n444), .A4(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(G113), .B(G122), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n477), .B(new_n356), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT90), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n439), .A2(G146), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n446), .ZN(new_n481));
  NAND2_X1  g295(.A1(KEYINPUT18), .A2(G131), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  AOI22_X1  g297(.A1(new_n479), .A2(new_n481), .B1(new_n470), .B2(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n468), .B(new_n482), .C1(new_n467), .C2(new_n469), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n480), .A2(KEYINPUT90), .A3(new_n446), .ZN(new_n486));
  AND2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  AND3_X1   g302(.A1(new_n476), .A2(new_n478), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT19), .ZN(new_n490));
  OAI211_X1 g304(.A(new_n429), .B(new_n430), .C1(KEYINPUT91), .C2(new_n490), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n429), .A2(new_n430), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n491), .B(new_n213), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n441), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n471), .A2(new_n473), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n496), .A2(new_n497), .B1(new_n484), .B2(new_n487), .ZN(new_n498));
  OR2_X1    g312(.A1(new_n498), .A2(KEYINPUT92), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n478), .B1(new_n498), .B2(KEYINPUT92), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n489), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(G475), .A2(G902), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT20), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n476), .A2(new_n478), .A3(new_n488), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n496), .A2(new_n497), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n506), .A2(KEYINPUT92), .A3(new_n488), .ZN(new_n507));
  INV_X1    g321(.A(new_n478), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n498), .A2(KEYINPUT92), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n505), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT20), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(new_n502), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n504), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT9), .B(G234), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n412), .A2(G953), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(KEYINPUT95), .B1(new_n209), .B2(G128), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT95), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(new_n211), .A3(G143), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n209), .A2(G128), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n226), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(G134), .A3(new_n521), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT13), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n520), .A2(new_n525), .A3(G134), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n523), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n520), .A2(new_n525), .A3(G134), .A4(new_n521), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n188), .A2(new_n190), .A3(G122), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT93), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n341), .A2(KEYINPUT93), .A3(G122), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n187), .A2(G122), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(G107), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n535), .A2(new_n352), .A3(new_n537), .ZN(new_n540));
  AOI21_X1  g354(.A(KEYINPUT94), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n352), .B1(new_n535), .B2(new_n537), .ZN(new_n542));
  AOI211_X1 g356(.A(G107), .B(new_n536), .C1(new_n533), .C2(new_n534), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT94), .ZN(new_n544));
  NOR3_X1   g358(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n530), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n536), .B1(new_n535), .B2(KEYINPUT14), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n547), .B1(KEYINPUT14), .B2(new_n535), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G107), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n523), .A2(new_n524), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n549), .A2(new_n540), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n516), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n539), .A2(KEYINPUT94), .A3(new_n540), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n544), .B1(new_n542), .B2(new_n543), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n529), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n540), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n548), .B2(G107), .ZN(new_n557));
  INV_X1    g371(.A(new_n516), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n323), .B1(new_n552), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(G478), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(KEYINPUT15), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n546), .A2(new_n551), .A3(new_n516), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n558), .B1(new_n555), .B2(new_n557), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n566), .B(new_n323), .C1(KEYINPUT15), .C2(new_n561), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n478), .B1(new_n476), .B2(new_n488), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n323), .B1(new_n489), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G475), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n514), .A2(new_n563), .A3(new_n567), .A4(new_n570), .ZN(new_n571));
  NOR4_X1   g385(.A1(new_n325), .A2(new_n410), .A3(new_n465), .A4(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(G221), .B1(new_n515), .B2(G902), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT85), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n367), .A2(new_n278), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(KEYINPUT84), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT84), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n367), .A2(new_n278), .A3(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n216), .B1(new_n223), .B2(new_n249), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n365), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n577), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n582), .A2(KEYINPUT12), .A3(new_n253), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT12), .B1(new_n582), .B2(new_n253), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n575), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT12), .ZN(new_n586));
  INV_X1    g400(.A(new_n579), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n580), .A2(new_n359), .A3(new_n364), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n578), .B1(new_n367), .B2(new_n278), .ZN(new_n589));
  NOR3_X1   g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n586), .B1(new_n590), .B2(new_n273), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n582), .A2(KEYINPUT12), .A3(new_n253), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n591), .A2(KEYINPUT85), .A3(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT10), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n581), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n381), .A2(new_n250), .A3(new_n383), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n365), .A2(KEYINPUT10), .A3(new_n224), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n253), .ZN(new_n599));
  XNOR2_X1  g413(.A(G110), .B(G140), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n449), .A2(G227), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n600), .B(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(KEYINPUT80), .B(KEYINPUT81), .ZN(new_n603));
  XOR2_X1   g417(.A(new_n602), .B(new_n603), .Z(new_n604));
  NOR2_X1   g418(.A1(new_n599), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n585), .A2(new_n593), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(KEYINPUT86), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT86), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n585), .A2(new_n593), .A3(new_n605), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n598), .B(new_n273), .ZN(new_n610));
  INV_X1    g424(.A(new_n604), .ZN(new_n611));
  OR2_X1    g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n607), .A2(new_n609), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(G469), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n613), .A2(new_n614), .A3(new_n323), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n610), .A2(new_n611), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n599), .B1(new_n591), .B2(new_n592), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n616), .B1(new_n611), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n614), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n614), .A2(new_n323), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n574), .B1(new_n615), .B2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n572), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(G101), .ZN(G3));
  OAI21_X1  g438(.A(G472), .B1(new_n291), .B2(G902), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n305), .A2(new_n292), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI211_X1 g441(.A(new_n574), .B(new_n627), .C1(new_n615), .C2(new_n621), .ZN(new_n628));
  INV_X1    g442(.A(new_n465), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n397), .A2(new_n406), .ZN(new_n631));
  INV_X1    g445(.A(new_n407), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n397), .A2(new_n406), .A3(new_n407), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n633), .A2(KEYINPUT96), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT96), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n336), .B1(new_n409), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n513), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n512), .B1(new_n511), .B2(new_n502), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n570), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n561), .A2(G902), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT97), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(KEYINPUT33), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n644), .A2(KEYINPUT33), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n566), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT33), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n564), .A2(new_n565), .A3(KEYINPUT97), .A4(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n643), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n560), .A2(new_n561), .ZN(new_n652));
  INV_X1    g466(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n641), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n638), .A2(new_n334), .A3(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n630), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT98), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT34), .B(G104), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G6));
  AND2_X1   g473(.A1(new_n635), .A2(new_n637), .ZN(new_n660));
  INV_X1    g474(.A(new_n641), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n563), .A2(new_n567), .ZN(new_n662));
  INV_X1    g476(.A(new_n334), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(KEYINPUT99), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n660), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT99), .B1(new_n638), .B2(new_n667), .ZN(new_n668));
  AND2_X1   g482(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n630), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT35), .B(G107), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G9));
  NOR2_X1   g487(.A1(new_n455), .A2(KEYINPUT36), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n448), .B(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n462), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n460), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n410), .A2(new_n571), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n628), .A2(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(KEYINPUT37), .B(G110), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G12));
  NOR2_X1   g496(.A1(new_n325), .A2(new_n678), .ZN(new_n683));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n332), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n329), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n661), .A2(new_n662), .A3(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n622), .A2(new_n683), .A3(new_n687), .A4(new_n660), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G128), .ZN(G30));
  XNOR2_X1  g503(.A(new_n686), .B(KEYINPUT39), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n622), .A2(new_n690), .ZN(new_n691));
  OR2_X1    g505(.A1(new_n691), .A2(KEYINPUT40), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(KEYINPUT40), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n408), .A2(new_n409), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(KEYINPUT38), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n633), .A2(new_n634), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT38), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n294), .A2(new_n307), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n262), .A2(new_n296), .ZN(new_n701));
  AOI22_X1  g515(.A1(new_n302), .A2(new_n268), .B1(new_n701), .B2(new_n290), .ZN(new_n702));
  OAI21_X1  g516(.A(G472), .B1(new_n702), .B2(G902), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  AOI22_X1  g518(.A1(new_n514), .A2(new_n570), .B1(new_n563), .B2(new_n567), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(new_n335), .A3(new_n678), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n699), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n692), .A2(new_n693), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT100), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G143), .ZN(G45));
  OAI211_X1 g524(.A(new_n641), .B(new_n686), .C1(new_n651), .C2(new_n653), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(KEYINPUT101), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n712), .A2(new_n622), .A3(new_n660), .A4(new_n683), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  AND3_X1   g528(.A1(new_n613), .A2(new_n614), .A3(new_n323), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n614), .B1(new_n613), .B2(new_n323), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n715), .A2(new_n716), .A3(new_n574), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n325), .A2(new_n465), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(new_n718), .A3(new_n655), .ZN(new_n719));
  XNOR2_X1  g533(.A(KEYINPUT41), .B(G113), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G15));
  NAND2_X1  g535(.A1(new_n717), .A2(new_n718), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n669), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(KEYINPUT102), .B(G116), .Z(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G18));
  NOR2_X1   g539(.A1(new_n571), .A2(new_n334), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n717), .A2(new_n660), .A3(new_n683), .A4(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G119), .ZN(G21));
  OAI21_X1  g542(.A(new_n311), .B1(new_n316), .B2(new_n317), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(new_n290), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n271), .A2(new_n272), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n292), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n734));
  INV_X1    g548(.A(new_n456), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n455), .B1(new_n442), .B2(new_n447), .ZN(new_n736));
  OAI21_X1  g550(.A(new_n323), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(new_n417), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n457), .A2(new_n323), .A3(new_n418), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n415), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n734), .B1(new_n740), .B2(new_n463), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n460), .A2(KEYINPUT103), .A3(new_n464), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AND4_X1   g557(.A1(new_n663), .A2(new_n733), .A3(new_n743), .A4(new_n625), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n635), .A2(new_n705), .A3(new_n637), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n613), .A2(new_n323), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(G469), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n573), .A3(new_n615), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n746), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n733), .A2(new_n743), .A3(new_n625), .A4(new_n663), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n635), .A2(new_n705), .A3(new_n637), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT104), .B1(new_n717), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n751), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(G122), .Z(G24));
  NAND2_X1  g571(.A1(new_n648), .A2(new_n650), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n642), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n652), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(KEYINPUT101), .A3(new_n641), .A4(new_n686), .ZN(new_n761));
  INV_X1    g575(.A(new_n678), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n733), .A2(new_n625), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT101), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n711), .A2(new_n764), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n761), .A2(new_n763), .A3(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n660), .A3(new_n717), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G125), .ZN(G27));
  INV_X1    g582(.A(KEYINPUT42), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n696), .A2(new_n336), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n573), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT106), .ZN(new_n772));
  OAI21_X1  g586(.A(KEYINPUT105), .B1(new_n617), .B2(new_n611), .ZN(new_n773));
  OAI22_X1  g587(.A1(new_n583), .A2(new_n584), .B1(new_n253), .B2(new_n598), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT105), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n775), .A3(new_n604), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n773), .A2(new_n776), .A3(G469), .A4(new_n616), .ZN(new_n777));
  INV_X1    g591(.A(new_n620), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n772), .B1(new_n715), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n779), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n615), .A3(KEYINPUT106), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n771), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n325), .ZN(new_n784));
  AND4_X1   g598(.A1(new_n784), .A2(new_n761), .A3(new_n765), .A4(new_n743), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n769), .B1(new_n783), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n771), .ZN(new_n787));
  AND3_X1   g601(.A1(new_n781), .A2(new_n615), .A3(KEYINPUT106), .ZN(new_n788));
  AOI21_X1  g602(.A(KEYINPUT106), .B1(new_n781), .B2(new_n615), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n718), .B(new_n787), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n712), .A2(new_n769), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT107), .B1(new_n786), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n784), .A2(new_n743), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n712), .A2(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n797));
  OAI21_X1  g611(.A(KEYINPUT42), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n783), .A2(new_n769), .A3(new_n718), .A4(new_n712), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT107), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n798), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n793), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(new_n230), .ZN(G33));
  NAND2_X1  g617(.A1(new_n780), .A2(new_n782), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n804), .A2(new_n718), .A3(new_n687), .A4(new_n787), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G134), .ZN(G36));
  INV_X1    g620(.A(KEYINPUT43), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n760), .A2(new_n807), .A3(new_n661), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n651), .A2(new_n653), .ZN(new_n809));
  OAI21_X1  g623(.A(KEYINPUT43), .B1(new_n809), .B2(new_n641), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n678), .B1(new_n625), .B2(new_n626), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT44), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n812), .A2(KEYINPUT44), .A3(new_n813), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n770), .A3(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT45), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n614), .B1(new_n618), .B2(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n773), .A2(new_n776), .A3(KEYINPUT45), .A4(new_n616), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n620), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n822), .A2(KEYINPUT46), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n615), .B1(new_n822), .B2(KEYINPUT46), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n825), .A2(new_n574), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(new_n690), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n818), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(KEYINPUT108), .B(G137), .Z(new_n829));
  XNOR2_X1  g643(.A(new_n828), .B(new_n829), .ZN(G39));
  NAND4_X1  g644(.A1(new_n712), .A2(new_n325), .A3(new_n465), .A4(new_n770), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT47), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n825), .B2(new_n574), .ZN(new_n833));
  OAI211_X1 g647(.A(KEYINPUT47), .B(new_n573), .C1(new_n823), .C2(new_n824), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(new_n428), .ZN(G42));
  AOI22_X1  g650(.A1(new_n628), .A2(new_n679), .B1(new_n572), .B2(new_n622), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT109), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n654), .A2(new_n838), .B1(new_n662), .B2(new_n661), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n760), .A2(KEYINPUT109), .A3(new_n641), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(new_n410), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n628), .A2(new_n841), .A3(new_n629), .A4(new_n842), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n837), .B(new_n843), .C1(new_n751), .C2(new_n755), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n719), .B(new_n727), .C1(new_n669), .C2(new_n722), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n783), .A2(new_n766), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n661), .A2(new_n563), .A3(new_n567), .A4(new_n686), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n694), .A2(new_n335), .ZN(new_n849));
  OR3_X1    g663(.A1(new_n848), .A2(new_n849), .A3(KEYINPUT110), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT110), .B1(new_n848), .B2(new_n849), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n850), .A2(new_n622), .A3(new_n683), .A4(new_n851), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n847), .A2(new_n805), .A3(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n846), .A2(new_n793), .A3(new_n801), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n678), .A2(new_n573), .A3(new_n686), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n704), .A2(new_n855), .ZN(new_n856));
  OAI211_X1 g670(.A(new_n856), .B(new_n745), .C1(new_n788), .C2(new_n789), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n767), .A2(new_n713), .A3(new_n857), .A4(new_n688), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT52), .ZN(new_n859));
  OAI21_X1  g673(.A(KEYINPUT53), .B1(new_n854), .B2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(new_n802), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT53), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n847), .A2(new_n805), .A3(new_n852), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n863), .A2(new_n844), .A3(new_n845), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n861), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n688), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n749), .A2(new_n638), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n866), .B1(new_n867), .B2(new_n766), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n868), .A2(KEYINPUT52), .A3(new_n713), .A4(new_n857), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT52), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n858), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n869), .A2(new_n871), .A3(KEYINPUT111), .ZN(new_n872));
  OR3_X1    g686(.A1(new_n858), .A2(KEYINPUT111), .A3(new_n870), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n860), .B(KEYINPUT54), .C1(new_n865), .C2(new_n874), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n715), .A2(new_n716), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n574), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n833), .A2(new_n834), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT112), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n733), .A2(new_n743), .A3(new_n625), .A4(new_n330), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n811), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n879), .B1(new_n881), .B2(new_n770), .ZN(new_n882));
  NOR4_X1   g696(.A1(new_n811), .A2(new_n849), .A3(new_n880), .A4(KEYINPUT112), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  NOR4_X1   g699(.A1(new_n771), .A2(new_n715), .A3(new_n329), .A4(new_n716), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n704), .A2(new_n629), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n661), .A3(new_n809), .A4(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n886), .A2(new_n763), .A3(new_n812), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n811), .A2(new_n880), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n699), .A2(new_n336), .ZN(new_n892));
  OAI21_X1  g706(.A(KEYINPUT113), .B1(new_n892), .B2(new_n749), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT113), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n717), .A2(new_n699), .A3(new_n894), .A4(new_n336), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n891), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(KEYINPUT50), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT50), .ZN(new_n898));
  AOI211_X1 g712(.A(new_n898), .B(new_n891), .C1(new_n893), .C2(new_n895), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n885), .B(new_n890), .C1(new_n897), .C2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(KEYINPUT51), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n896), .B(KEYINPUT50), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(KEYINPUT51), .A3(new_n885), .A4(new_n890), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n886), .A2(new_n795), .A3(new_n812), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT114), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n906), .A2(KEYINPUT48), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(KEYINPUT48), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n905), .B2(new_n908), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n867), .A2(new_n881), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n886), .A2(new_n887), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n327), .B(new_n911), .C1(new_n912), .C2(new_n654), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  AND3_X1   g728(.A1(new_n902), .A2(new_n904), .A3(new_n914), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n862), .B1(new_n854), .B2(new_n859), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n786), .A2(new_n792), .A3(new_n862), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n872), .A2(new_n873), .A3(new_n864), .A4(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n875), .A2(new_n915), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n326), .A2(new_n449), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI211_X1 g737(.A(new_n574), .B(new_n336), .C1(new_n741), .C2(new_n742), .ZN(new_n924));
  AND4_X1   g738(.A1(new_n661), .A2(new_n704), .A3(new_n760), .A4(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT49), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n876), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT49), .B1(new_n715), .B2(new_n716), .ZN(new_n928));
  NAND4_X1  g742(.A1(new_n925), .A2(new_n699), .A3(new_n927), .A4(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n923), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(KEYINPUT115), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT115), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n923), .A2(new_n932), .A3(new_n929), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(G75));
  NOR2_X1   g748(.A1(new_n449), .A2(G952), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT118), .Z(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n916), .A2(new_n919), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n938), .A2(new_n264), .A3(new_n323), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n401), .A2(new_n403), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT116), .Z(new_n941));
  XNOR2_X1  g755(.A(new_n405), .B(KEYINPUT117), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT55), .Z(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(new_n944), .ZN(new_n945));
  OR3_X1    g759(.A1(new_n939), .A2(KEYINPUT56), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n945), .B1(new_n939), .B2(KEYINPUT56), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n937), .B1(new_n946), .B2(new_n947), .ZN(G51));
  XNOR2_X1  g762(.A(new_n620), .B(KEYINPUT57), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n916), .A2(new_n917), .A3(new_n919), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n917), .B1(new_n916), .B2(new_n919), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT119), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI211_X1 g768(.A(KEYINPUT119), .B(new_n949), .C1(new_n950), .C2(new_n951), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n613), .A3(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n938), .A2(new_n323), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n957), .A2(new_n821), .A3(new_n820), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n935), .B1(new_n956), .B2(new_n958), .ZN(G54));
  NAND3_X1  g773(.A1(new_n957), .A2(KEYINPUT58), .A3(G475), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n960), .A2(new_n501), .ZN(new_n961));
  INV_X1    g775(.A(new_n935), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n957), .A2(KEYINPUT58), .A3(G475), .A4(new_n511), .ZN(new_n963));
  AND3_X1   g777(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(G60));
  XOR2_X1   g778(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n965));
  NOR2_X1   g779(.A1(new_n561), .A2(new_n323), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n758), .B(new_n967), .C1(new_n950), .C2(new_n951), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(new_n936), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n875), .A2(new_n920), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n758), .B1(new_n970), .B2(new_n967), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n969), .A2(new_n971), .ZN(G63));
  XNOR2_X1  g786(.A(KEYINPUT121), .B(KEYINPUT60), .ZN(new_n973));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n461), .B1(new_n938), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n975), .B1(new_n916), .B2(new_n919), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n937), .B1(new_n977), .B2(new_n675), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n978), .A2(KEYINPUT122), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n979), .A2(new_n980), .A3(KEYINPUT61), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n976), .B(new_n978), .C1(KEYINPUT122), .C2(new_n982), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n981), .A2(new_n983), .ZN(G66));
  OAI21_X1  g798(.A(G953), .B1(new_n333), .B2(new_n389), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n846), .B(KEYINPUT123), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n985), .B1(new_n987), .B2(G953), .ZN(new_n988));
  INV_X1    g802(.A(new_n941), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n989), .B1(G898), .B2(new_n449), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n988), .B(new_n990), .ZN(G69));
  OAI21_X1  g805(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n992), .B(KEYINPUT124), .Z(new_n993));
  XOR2_X1   g807(.A(new_n301), .B(new_n993), .Z(new_n994));
  INV_X1    g808(.A(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n868), .A2(new_n713), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT125), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n709), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(KEYINPUT62), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT62), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n997), .A2(new_n1000), .A3(new_n709), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n841), .A2(new_n718), .A3(new_n770), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n828), .B1(new_n691), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n1003), .A2(new_n835), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n999), .A2(new_n1001), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n995), .B1(new_n1005), .B2(new_n449), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n449), .B1(G227), .B2(G900), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT126), .Z(new_n1008));
  NAND4_X1  g822(.A1(new_n826), .A2(new_n690), .A3(new_n745), .A4(new_n795), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n1009), .B(new_n805), .C1(new_n818), .C2(new_n827), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n1010), .A2(new_n835), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n997), .A2(new_n1011), .A3(new_n861), .ZN(new_n1012));
  NAND2_X1  g826(.A1(new_n1012), .A2(new_n449), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n684), .A2(G953), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n994), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OR3_X1    g829(.A1(new_n1006), .A2(new_n1008), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1008), .B1(new_n1006), .B2(new_n1015), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(G72));
  NAND2_X1  g832(.A1(G472), .A2(G902), .ZN(new_n1019));
  XOR2_X1   g833(.A(new_n1019), .B(KEYINPUT63), .Z(new_n1020));
  OAI21_X1  g834(.A(new_n1020), .B1(new_n1012), .B2(new_n986), .ZN(new_n1021));
  NOR3_X1   g835(.A1(new_n320), .A2(new_n282), .A3(new_n268), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n935), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n860), .B1(new_n865), .B2(new_n874), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n321), .A2(new_n269), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1025), .A2(new_n1020), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1023), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1027));
  NAND4_X1  g841(.A1(new_n999), .A2(new_n987), .A3(new_n1004), .A4(new_n1001), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n1020), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n302), .A2(new_n312), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1031), .A2(KEYINPUT127), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT127), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1029), .A2(new_n1033), .A3(new_n1030), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1027), .B1(new_n1032), .B2(new_n1034), .ZN(G57));
endmodule


