//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n207));
  INV_X1    g0007(.A(G226), .ZN(new_n208));
  INV_X1    g0008(.A(G87), .ZN(new_n209));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  OAI221_X1 g0010(.A(new_n207), .B1(new_n202), .B2(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n206), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(KEYINPUT1), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n206), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XOR2_X1   g0019(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n220));
  XNOR2_X1  g0020(.A(new_n219), .B(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  INV_X1    g0022(.A(G20), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n201), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(G50), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n221), .B1(new_n225), .B2(new_n227), .C1(KEYINPUT1), .C2(new_n215), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n217), .A2(new_n228), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G250), .B(G257), .Z(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G116), .Z(new_n238));
  XNOR2_X1  g0038(.A(G97), .B(G107), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n202), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n240), .B(new_n246), .ZN(G351));
  XNOR2_X1  g0047(.A(KEYINPUT3), .B(G33), .ZN(new_n248));
  INV_X1    g0048(.A(G1698), .ZN(new_n249));
  NAND3_X1  g0049(.A1(new_n248), .A2(G222), .A3(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n248), .A2(G223), .A3(G1698), .ZN(new_n251));
  INV_X1    g0051(.A(G77), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n250), .B(new_n251), .C1(new_n252), .C2(new_n248), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(KEYINPUT66), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT66), .ZN(new_n257));
  NAND4_X1  g0057(.A1(new_n254), .A2(new_n257), .A3(G1), .A4(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n253), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n261), .B(G274), .C1(G41), .C2(G45), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n261), .B1(G41), .B2(G45), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n255), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n262), .B1(new_n264), .B2(new_n208), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n260), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G190), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT9), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n203), .A2(G20), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT67), .ZN(new_n271));
  XOR2_X1   g0071(.A(KEYINPUT8), .B(G58), .Z(new_n272));
  INV_X1    g0072(.A(G33), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(G20), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT67), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n203), .A2(new_n276), .A3(G20), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G20), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G150), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n271), .A2(new_n275), .A3(new_n277), .A4(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(new_n222), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n223), .A2(G1), .ZN(new_n284));
  NOR3_X1   g0084(.A1(new_n282), .A2(new_n284), .A3(new_n202), .ZN(new_n285));
  NAND3_X1  g0085(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n285), .B1(new_n202), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n283), .A2(new_n288), .ZN(new_n289));
  OAI22_X1  g0089(.A1(new_n267), .A2(new_n268), .B1(new_n269), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n289), .A2(new_n269), .ZN(new_n291));
  INV_X1    g0091(.A(G200), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n291), .B1(new_n292), .B2(new_n266), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT10), .B1(new_n290), .B2(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n289), .ZN(new_n295));
  AOI22_X1  g0095(.A1(KEYINPUT9), .A2(new_n295), .B1(new_n266), .B2(G190), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n267), .A2(G200), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n296), .A2(new_n297), .A3(new_n298), .A4(new_n291), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n272), .A2(new_n278), .B1(G20), .B2(G77), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n223), .A2(G33), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT15), .B(G87), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n284), .A2(KEYINPUT69), .A3(G13), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT69), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n286), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  AOI22_X1  g0108(.A1(new_n304), .A2(new_n282), .B1(new_n252), .B2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n282), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n305), .A2(new_n310), .A3(new_n307), .ZN(new_n311));
  INV_X1    g0111(.A(new_n284), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(G77), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n309), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(G244), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n262), .B1(new_n264), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n248), .A2(G232), .A3(new_n249), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n248), .A2(G238), .A3(G1698), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n273), .A2(KEYINPUT3), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT3), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n320), .A2(G33), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G107), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n317), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  OR2_X1    g0124(.A1(new_n324), .A2(KEYINPUT68), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n324), .A2(KEYINPUT68), .B1(new_n256), .B2(new_n258), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n316), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n314), .B1(new_n327), .B2(G190), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n327), .A2(new_n292), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G179), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n266), .A2(new_n331), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n332), .B(new_n289), .C1(G169), .C2(new_n266), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n300), .A2(new_n330), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT7), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n248), .A2(new_n335), .A3(G20), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT7), .B1(new_n322), .B2(new_n223), .ZN(new_n337));
  OAI21_X1  g0137(.A(G68), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G58), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(new_n242), .ZN(new_n340));
  OAI21_X1  g0140(.A(G20), .B1(new_n340), .B2(new_n201), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n278), .A2(G159), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n338), .A2(KEYINPUT16), .A3(new_n344), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT16), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n335), .B1(new_n248), .B2(G20), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n322), .A2(KEYINPUT7), .A3(new_n223), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n242), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n346), .B1(new_n349), .B2(new_n343), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n345), .A2(new_n350), .A3(new_n282), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT8), .B(G58), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n352), .A2(new_n282), .A3(new_n284), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(new_n287), .B2(new_n352), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(G232), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n262), .B1(new_n264), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT74), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n319), .A2(new_n321), .A3(G226), .A4(G1698), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n319), .A2(new_n321), .A3(G223), .A4(new_n249), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G87), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n259), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT74), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n364), .B(new_n262), .C1(new_n264), .C2(new_n356), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n358), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n357), .B1(new_n259), .B2(new_n362), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(G169), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n366), .A2(new_n331), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n355), .A2(KEYINPUT18), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g0172(.A(KEYINPUT18), .B1(new_n355), .B2(new_n370), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n358), .A2(new_n363), .A3(new_n365), .ZN(new_n375));
  OAI22_X1  g0175(.A1(new_n375), .A2(G190), .B1(G200), .B2(new_n367), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n376), .A2(new_n351), .A3(new_n354), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT17), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n377), .B(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n314), .B1(new_n327), .B2(G169), .ZN(new_n380));
  AOI21_X1  g0180(.A(KEYINPUT70), .B1(new_n327), .B2(new_n331), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n327), .A2(KEYINPUT70), .A3(new_n331), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n380), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NOR4_X1   g0184(.A1(new_n334), .A2(new_n374), .A3(new_n379), .A4(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT12), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n386), .A2(G68), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n308), .A2(new_n387), .B1(new_n386), .B2(new_n286), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n386), .B1(new_n311), .B2(new_n312), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT11), .ZN(new_n390));
  AOI22_X1  g0190(.A1(new_n274), .A2(G77), .B1(G20), .B2(new_n242), .ZN(new_n391));
  INV_X1    g0191(.A(new_n278), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n391), .B1(new_n202), .B2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n390), .B1(new_n393), .B2(new_n282), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n393), .A2(new_n390), .A3(new_n282), .ZN(new_n395));
  OAI221_X1 g0195(.A(new_n388), .B1(new_n389), .B2(new_n242), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n255), .A2(G238), .A3(new_n263), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n262), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT71), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n397), .A2(KEYINPUT71), .A3(new_n262), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT13), .ZN(new_n403));
  NOR3_X1   g0203(.A1(new_n322), .A2(new_n356), .A3(new_n249), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n319), .A2(new_n321), .A3(G226), .A4(new_n249), .ZN(new_n405));
  NAND2_X1  g0205(.A1(G33), .A2(G97), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n259), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  AND3_X1   g0208(.A1(new_n402), .A2(new_n403), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n403), .B1(new_n402), .B2(new_n408), .ZN(new_n410));
  OAI21_X1  g0210(.A(G169), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(KEYINPUT14), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT14), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n413), .B(G169), .C1(new_n409), .C2(new_n410), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n402), .A2(new_n408), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(KEYINPUT13), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT72), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n402), .A2(new_n403), .A3(new_n408), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n402), .A2(KEYINPUT72), .A3(new_n403), .A4(new_n408), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n331), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n396), .B1(new_n415), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(new_n421), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G190), .ZN(new_n425));
  OAI21_X1  g0225(.A(G200), .B1(new_n409), .B2(new_n410), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n388), .B1(new_n395), .B2(new_n394), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n311), .A2(new_n312), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n242), .B1(new_n428), .B2(KEYINPUT12), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n431), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT73), .B1(new_n425), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n268), .B1(new_n420), .B2(new_n421), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT73), .ZN(new_n435));
  NOR3_X1   g0235(.A1(new_n434), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n423), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n385), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g0239(.A(KEYINPUT5), .B(G41), .ZN(new_n440));
  INV_X1    g0240(.A(G45), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(G1), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(G274), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n445), .B1(new_n442), .B2(new_n440), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n446), .B2(G270), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n319), .A2(new_n321), .A3(G257), .A4(new_n249), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n319), .A2(new_n321), .A3(G264), .A4(G1698), .ZN(new_n449));
  INV_X1    g0249(.A(G303), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n448), .B(new_n449), .C1(new_n450), .C2(new_n248), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n451), .A2(KEYINPUT79), .A3(new_n259), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT79), .B1(new_n451), .B2(new_n259), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n447), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G116), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n308), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g0256(.A(new_n455), .B1(new_n261), .B2(G33), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n305), .A2(new_n310), .A3(new_n307), .A4(new_n457), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G283), .ZN(new_n460));
  INV_X1    g0260(.A(G97), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n460), .B(new_n223), .C1(G33), .C2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n455), .A2(G20), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n282), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT20), .ZN(new_n465));
  XNOR2_X1  g0265(.A(new_n464), .B(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n369), .B1(new_n459), .B2(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n454), .A2(new_n467), .A3(KEYINPUT21), .ZN(new_n468));
  AOI21_X1  g0268(.A(KEYINPUT21), .B1(new_n454), .B2(new_n467), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n446), .A2(G270), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n443), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n451), .A2(new_n259), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT79), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n451), .A2(KEYINPUT79), .A3(new_n259), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AND2_X1   g0277(.A1(new_n464), .A2(new_n465), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n464), .A2(new_n465), .ZN(new_n479));
  OAI211_X1 g0279(.A(new_n458), .B(new_n456), .C1(new_n478), .C2(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n477), .A2(KEYINPUT80), .A3(G179), .A4(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT80), .ZN(new_n482));
  OAI211_X1 g0282(.A(G179), .B(new_n447), .C1(new_n452), .C2(new_n453), .ZN(new_n483));
  INV_X1    g0283(.A(new_n480), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n454), .A2(G200), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n486), .B(new_n484), .C1(new_n268), .C2(new_n454), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n470), .A2(new_n481), .A3(new_n485), .A4(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n261), .A2(G33), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n286), .A2(new_n489), .A3(new_n222), .A4(new_n281), .ZN(new_n490));
  AND2_X1   g0290(.A1(new_n490), .A2(KEYINPUT75), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n490), .A2(KEYINPUT75), .ZN(new_n492));
  OAI21_X1  g0292(.A(G87), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT19), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n223), .B1(new_n406), .B2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(G107), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n209), .A2(new_n461), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n319), .A2(new_n321), .A3(new_n223), .A4(G68), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n494), .B1(new_n302), .B2(new_n461), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n501), .A2(new_n282), .B1(new_n308), .B2(new_n303), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n442), .A2(G274), .ZN(new_n504));
  OAI21_X1  g0304(.A(G250), .B1(new_n441), .B2(G1), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n504), .B1(new_n445), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g0306(.A1(new_n319), .A2(new_n321), .A3(G244), .A4(G1698), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n319), .A2(new_n321), .A3(G238), .A4(new_n249), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G116), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n506), .B1(new_n510), .B2(new_n259), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n511), .A2(new_n292), .ZN(new_n512));
  AOI211_X1 g0312(.A(new_n268), .B(new_n506), .C1(new_n510), .C2(new_n259), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n503), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n510), .A2(new_n259), .ZN(new_n515));
  INV_X1    g0315(.A(new_n506), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G169), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n511), .A2(G179), .ZN(new_n519));
  INV_X1    g0319(.A(new_n303), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n491), .B2(new_n492), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n518), .A2(new_n519), .B1(new_n521), .B2(new_n502), .ZN(new_n522));
  OAI21_X1  g0322(.A(KEYINPUT78), .B1(new_n514), .B2(new_n522), .ZN(new_n523));
  OAI21_X1  g0323(.A(G107), .B1(new_n491), .B2(new_n492), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT81), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT25), .ZN(new_n526));
  AOI21_X1  g0326(.A(G107), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n287), .B(new_n527), .C1(new_n525), .C2(new_n526), .ZN(new_n528));
  OAI211_X1 g0328(.A(KEYINPUT81), .B(KEYINPUT25), .C1(new_n286), .C2(G107), .ZN(new_n529));
  AND2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n524), .A2(new_n530), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n319), .A2(new_n321), .A3(new_n223), .A4(G87), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n532), .A2(KEYINPUT22), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT22), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n248), .A2(new_n534), .A3(new_n223), .A4(G87), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT23), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n223), .B2(G107), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n496), .A2(KEYINPUT23), .A3(G20), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(G20), .B2(new_n509), .ZN(new_n541));
  INV_X1    g0341(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT24), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n310), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n541), .B1(new_n533), .B2(new_n535), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(KEYINPUT24), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n531), .B1(new_n545), .B2(new_n547), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n319), .A2(new_n321), .A3(G250), .A4(new_n249), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n319), .A2(new_n321), .A3(G257), .A4(G1698), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G294), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(new_n259), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n446), .A2(G264), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n553), .A2(new_n554), .A3(new_n443), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT82), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n556), .A3(new_n292), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(G190), .B2(new_n555), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n556), .B1(new_n555), .B2(new_n292), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n548), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n517), .A2(G200), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n511), .A2(G190), .ZN(new_n562));
  NAND4_X1  g0362(.A1(new_n561), .A2(new_n502), .A3(new_n493), .A4(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT78), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n521), .A2(new_n502), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n511), .A2(new_n369), .ZN(new_n566));
  AOI211_X1 g0366(.A(new_n331), .B(new_n506), .C1(new_n510), .C2(new_n259), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n282), .B1(new_n546), .B2(KEYINPUT24), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n543), .A2(new_n544), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n524), .B(new_n530), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n555), .A2(new_n369), .ZN(new_n573));
  AOI22_X1  g0373(.A1(new_n259), .A2(new_n552), .B1(new_n446), .B2(G264), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(new_n331), .A3(new_n443), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n523), .A2(new_n560), .A3(new_n569), .A4(new_n576), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n488), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n319), .A2(new_n321), .A3(G244), .A4(new_n249), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT4), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n248), .A2(KEYINPUT4), .A3(G244), .A4(new_n249), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n248), .A2(G250), .A3(G1698), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n460), .A4(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n259), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n444), .B1(new_n446), .B2(G257), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n369), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n440), .A2(new_n442), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n589), .A2(G257), .A3(new_n255), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n443), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n259), .B2(new_n584), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n331), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT6), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n594), .A2(new_n461), .A3(G107), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n595), .B1(new_n594), .B2(new_n239), .ZN(new_n596));
  OAI22_X1  g0396(.A1(new_n596), .A2(new_n223), .B1(new_n252), .B2(new_n392), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n496), .B1(new_n347), .B2(new_n348), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n282), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n286), .A2(G97), .ZN(new_n600));
  XNOR2_X1  g0400(.A(new_n490), .B(KEYINPUT75), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n600), .B1(new_n601), .B2(G97), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n588), .A2(new_n593), .A3(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT76), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n585), .A2(G190), .A3(new_n586), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(new_n599), .A3(new_n602), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n592), .A2(new_n292), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n605), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n599), .A2(new_n602), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n587), .A2(G200), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n610), .A2(new_n611), .A3(KEYINPUT76), .A4(new_n606), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n604), .B1(new_n609), .B2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT77), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI211_X1 g0415(.A(KEYINPUT77), .B(new_n604), .C1(new_n609), .C2(new_n612), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n578), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n439), .A2(new_n617), .ZN(G372));
  INV_X1    g0418(.A(new_n333), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n355), .A2(new_n370), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT18), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n371), .ZN(new_n623));
  INV_X1    g0423(.A(new_n423), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n425), .A2(new_n432), .A3(KEYINPUT73), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n435), .B1(new_n434), .B2(new_n431), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n624), .B1(new_n627), .B2(new_n384), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n623), .B1(new_n628), .B2(new_n379), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n619), .B1(new_n629), .B2(new_n300), .ZN(new_n630));
  OAI21_X1  g0430(.A(KEYINPUT83), .B1(new_n566), .B2(new_n567), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT83), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n519), .B(new_n632), .C1(new_n369), .C2(new_n511), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n631), .A2(new_n633), .B1(new_n521), .B2(new_n502), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n588), .A2(new_n593), .A3(new_n603), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n634), .A2(new_n635), .A3(new_n514), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n634), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n523), .A2(new_n604), .A3(new_n569), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n454), .A2(new_n467), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT21), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n454), .A2(new_n467), .A3(KEYINPUT21), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n643), .A2(new_n485), .A3(new_n481), .A4(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n576), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n609), .A2(new_n612), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n631), .A2(new_n633), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n514), .B1(new_n649), .B2(new_n565), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n648), .A2(new_n635), .A3(new_n560), .A4(new_n650), .ZN(new_n651));
  OAI211_X1 g0451(.A(new_n638), .B(new_n640), .C1(new_n647), .C2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n630), .B1(new_n439), .B2(new_n653), .ZN(G369));
  NAND3_X1  g0454(.A1(new_n261), .A2(new_n223), .A3(G13), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(KEYINPUT27), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT84), .ZN(new_n657));
  OAI21_X1  g0457(.A(G213), .B1(new_n655), .B2(KEYINPUT27), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G343), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n560), .B(new_n576), .C1(new_n548), .C2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n660), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n646), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n484), .A2(new_n660), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n645), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n488), .B2(new_n665), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G330), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n668), .A2(KEYINPUT85), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT85), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n671), .B1(new_n667), .B2(G330), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n664), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n645), .A2(new_n660), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n560), .A2(new_n576), .ZN(new_n676));
  XNOR2_X1  g0476(.A(new_n660), .B(KEYINPUT86), .ZN(new_n677));
  OAI22_X1  g0477(.A1(new_n675), .A2(new_n676), .B1(new_n576), .B2(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n674), .A2(new_n678), .ZN(G399));
  INV_X1    g0479(.A(new_n218), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(G41), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n497), .A2(G116), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(G1), .A3(new_n683), .ZN(new_n684));
  OAI21_X1  g0484(.A(new_n684), .B1(new_n227), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g0485(.A(new_n685), .B(KEYINPUT28), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT29), .ZN(new_n687));
  INV_X1    g0487(.A(new_n677), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n652), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  OAI21_X1  g0489(.A(KEYINPUT90), .B1(new_n651), .B2(new_n647), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n649), .A2(new_n565), .ZN(new_n691));
  AND2_X1   g0491(.A1(new_n650), .A2(new_n560), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n470), .A2(new_n481), .A3(new_n485), .A4(new_n576), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT90), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n692), .A2(new_n693), .A3(new_n694), .A4(new_n613), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n690), .A2(new_n691), .A3(new_n695), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n639), .A2(KEYINPUT89), .A3(new_n637), .ZN(new_n697));
  AOI21_X1  g0497(.A(KEYINPUT89), .B1(new_n639), .B2(new_n637), .ZN(new_n698));
  NOR4_X1   g0498(.A1(new_n634), .A2(new_n635), .A3(new_n637), .A4(new_n514), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n697), .A2(new_n698), .A3(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n660), .B1(new_n696), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n689), .B1(new_n701), .B2(KEYINPUT29), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n585), .A2(new_n574), .A3(new_n586), .A4(new_n511), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n703), .B1(new_n483), .B2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(KEYINPUT88), .ZN(new_n706));
  OR3_X1    g0506(.A1(new_n483), .A2(new_n704), .A3(new_n703), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT88), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n708), .B(new_n703), .C1(new_n483), .C2(new_n704), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n511), .A2(G179), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n454), .A2(new_n710), .A3(new_n587), .A4(new_n555), .ZN(new_n711));
  NAND4_X1  g0511(.A1(new_n706), .A2(new_n707), .A3(new_n709), .A4(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(KEYINPUT31), .B1(new_n712), .B2(new_n662), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n707), .A2(new_n705), .A3(new_n711), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n677), .A2(KEYINPUT31), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n714), .A2(new_n715), .A3(KEYINPUT87), .ZN(new_n716));
  AOI21_X1  g0516(.A(KEYINPUT87), .B1(new_n714), .B2(new_n715), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n713), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n578), .B(new_n688), .C1(new_n615), .C2(new_n616), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n669), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  AND2_X1   g0521(.A1(new_n702), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n686), .B1(new_n722), .B2(G1), .ZN(G364));
  NOR2_X1   g0523(.A1(new_n670), .A2(new_n672), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n223), .A2(G13), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n261), .B1(new_n725), .B2(G45), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n681), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  OAI211_X1 g0529(.A(new_n724), .B(new_n729), .C1(G330), .C2(new_n667), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n680), .A2(new_n322), .ZN(new_n731));
  AOI22_X1  g0531(.A1(new_n731), .A2(G355), .B1(new_n455), .B2(new_n680), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n322), .A2(new_n218), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT91), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(G45), .B2(new_n227), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n246), .A2(new_n441), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n732), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT92), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n222), .B1(G20), .B2(new_n369), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n729), .B1(new_n737), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g0545(.A(new_n745), .B(KEYINPUT93), .ZN(new_n746));
  INV_X1    g0546(.A(new_n743), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n223), .A2(G190), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G179), .A2(G200), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G329), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n322), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n331), .A2(new_n292), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n223), .A2(new_n268), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(G326), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n292), .A2(G179), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n755), .A2(new_n756), .B1(new_n758), .B2(new_n450), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n223), .B1(new_n749), .B2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI211_X1 g0561(.A(new_n752), .B(new_n759), .C1(G294), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n753), .A2(new_n748), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  XNOR2_X1  g0564(.A(KEYINPUT33), .B(G317), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n748), .A2(new_n757), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n764), .A2(new_n765), .B1(new_n767), .B2(G283), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n331), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n754), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n748), .A2(new_n769), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G322), .A2(new_n771), .B1(new_n773), .B2(G311), .ZN(new_n774));
  NAND3_X1  g0574(.A1(new_n762), .A2(new_n768), .A3(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(KEYINPUT94), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n755), .ZN(new_n778));
  AOI22_X1  g0578(.A1(G50), .A2(new_n778), .B1(new_n771), .B2(G58), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n252), .B2(new_n772), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n248), .B1(new_n758), .B2(new_n209), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n763), .A2(new_n242), .B1(new_n766), .B2(new_n496), .ZN(new_n782));
  NOR3_X1   g0582(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g0583(.A(G159), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n750), .A2(KEYINPUT32), .A3(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(KEYINPUT32), .ZN(new_n786));
  INV_X1    g0586(.A(new_n750), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n786), .B1(new_n787), .B2(G159), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n785), .B(new_n788), .C1(G97), .C2(new_n761), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n775), .A2(new_n776), .B1(new_n783), .B2(new_n789), .ZN(new_n790));
  AND2_X1   g0590(.A1(new_n777), .A2(new_n790), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n746), .B1(new_n747), .B2(new_n791), .C1(new_n667), .C2(new_n741), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n730), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(G396));
  INV_X1    g0594(.A(KEYINPUT98), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n651), .A2(new_n647), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n650), .A2(new_n637), .A3(new_n604), .ZN(new_n797));
  AND3_X1   g0597(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n564), .B1(new_n563), .B2(new_n568), .ZN(new_n799));
  NOR3_X1   g0599(.A1(new_n798), .A2(new_n799), .A3(new_n635), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n691), .B(new_n797), .C1(new_n800), .C2(new_n637), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n688), .B1(new_n796), .B2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n380), .ZN(new_n803));
  INV_X1    g0603(.A(new_n383), .ZN(new_n804));
  OAI211_X1 g0604(.A(new_n803), .B(new_n660), .C1(new_n804), .C2(new_n381), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n328), .A2(new_n329), .B1(new_n314), .B2(new_n662), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n805), .B1(new_n384), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n807), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n809), .B(new_n688), .C1(new_n796), .C2(new_n801), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n795), .B1(new_n721), .B2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n728), .B1(new_n721), .B2(new_n811), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n720), .A2(KEYINPUT98), .A3(new_n808), .A4(new_n810), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT99), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n747), .A2(new_n739), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n728), .B1(new_n817), .B2(G77), .ZN(new_n818));
  INV_X1    g0618(.A(G294), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n770), .A2(new_n819), .B1(new_n760), .B2(new_n461), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(KEYINPUT95), .Z(new_n821));
  INV_X1    g0621(.A(G283), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n755), .A2(new_n450), .B1(new_n763), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n758), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(G107), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n248), .B1(new_n773), .B2(G116), .ZN(new_n826));
  AOI22_X1  g0626(.A1(G87), .A2(new_n767), .B1(new_n787), .B2(G311), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n821), .A2(new_n825), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(G143), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n770), .A2(new_n829), .B1(new_n772), .B2(new_n784), .ZN(new_n830));
  AOI22_X1  g0630(.A1(G137), .A2(new_n778), .B1(new_n764), .B2(G150), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n831), .A2(KEYINPUT96), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(KEYINPUT96), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  XOR2_X1   g0634(.A(KEYINPUT97), .B(KEYINPUT34), .Z(new_n835));
  AND2_X1   g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(G132), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n248), .B1(new_n750), .B2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n767), .A2(G68), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n202), .B2(new_n758), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n838), .B(new_n840), .C1(G58), .C2(new_n761), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n834), .B2(new_n835), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n828), .B1(new_n836), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n818), .B1(new_n843), .B2(new_n743), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n809), .B2(new_n739), .ZN(new_n845));
  AND3_X1   g0645(.A1(new_n815), .A2(new_n816), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n816), .B1(new_n815), .B2(new_n845), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G384));
  INV_X1    g0649(.A(new_n596), .ZN(new_n850));
  OAI211_X1 g0650(.A(G116), .B(new_n224), .C1(new_n850), .C2(KEYINPUT35), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n851), .B1(KEYINPUT35), .B2(new_n850), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n852), .B(KEYINPUT36), .ZN(new_n853));
  OR3_X1    g0653(.A1(new_n227), .A2(new_n252), .A3(new_n340), .ZN(new_n854));
  AOI211_X1 g0654(.A(new_n261), .B(G13), .C1(new_n854), .C2(new_n241), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n355), .A2(KEYINPUT100), .A3(new_n370), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT100), .B1(new_n355), .B2(new_n370), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(new_n659), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n861), .B1(new_n351), .B2(new_n354), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  XOR2_X1   g0663(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n863), .A2(new_n377), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n863), .A2(new_n620), .A3(new_n377), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n860), .A2(new_n866), .B1(KEYINPUT37), .B2(new_n867), .ZN(new_n868));
  XNOR2_X1  g0668(.A(new_n377), .B(KEYINPUT17), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n863), .B1(new_n869), .B2(new_n623), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT38), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n862), .B1(new_n374), .B2(new_n379), .ZN(new_n873));
  INV_X1    g0673(.A(new_n355), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n862), .B1(new_n874), .B2(new_n376), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT100), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n620), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n875), .A2(new_n877), .A3(new_n865), .A4(new_n857), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n867), .A2(KEYINPUT37), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT38), .B1(new_n873), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT39), .B1(new_n872), .B2(new_n881), .ZN(new_n882));
  AOI22_X1  g0682(.A1(new_n860), .A2(new_n866), .B1(new_n867), .B2(new_n864), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n871), .B1(new_n883), .B2(new_n870), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n873), .A2(new_n880), .A3(KEYINPUT38), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT39), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n882), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n423), .A2(new_n662), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n430), .A2(new_n660), .ZN(new_n891));
  INV_X1    g0691(.A(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n627), .A2(new_n423), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n437), .A2(new_n891), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n810), .A2(new_n805), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n871), .B1(new_n868), .B2(new_n870), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n885), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n374), .A2(new_n861), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n890), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  XOR2_X1   g0700(.A(new_n900), .B(KEYINPUT104), .Z(new_n901));
  OAI21_X1  g0701(.A(new_n630), .B1(new_n702), .B2(new_n439), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n901), .B(new_n902), .ZN(new_n903));
  OR2_X1    g0703(.A1(KEYINPUT103), .A2(KEYINPUT31), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n712), .A2(new_n662), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n904), .B1(new_n712), .B2(new_n662), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n719), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n894), .A2(new_n893), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n897), .A2(new_n908), .A3(new_n909), .A4(new_n809), .ZN(new_n910));
  XOR2_X1   g0710(.A(KEYINPUT102), .B(KEYINPUT40), .Z(new_n911));
  NAND2_X1  g0711(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n913), .B1(new_n884), .B2(new_n885), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n914), .A2(new_n809), .A3(new_n909), .A4(new_n908), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n912), .A2(new_n915), .A3(G330), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n908), .A2(new_n385), .A3(G330), .A4(new_n438), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n908), .A2(new_n909), .A3(new_n809), .ZN(new_n918));
  AOI22_X1  g0718(.A1(new_n918), .A2(new_n914), .B1(new_n910), .B2(new_n911), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n439), .B1(new_n719), .B2(new_n907), .ZN(new_n920));
  AOI22_X1  g0720(.A1(new_n916), .A2(new_n917), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n903), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n922), .B1(new_n261), .B2(new_n725), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n903), .A2(new_n921), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n856), .B1(new_n923), .B2(new_n924), .ZN(G367));
  OAI21_X1  g0725(.A(new_n613), .B1(new_n610), .B2(new_n688), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n604), .A2(new_n677), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n675), .A2(new_n676), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT42), .Z(new_n931));
  OAI21_X1  g0731(.A(new_n635), .B1(new_n926), .B2(new_n576), .ZN(new_n932));
  AND2_X1   g0732(.A1(new_n932), .A2(KEYINPUT105), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n932), .A2(KEYINPUT105), .ZN(new_n934));
  NOR3_X1   g0734(.A1(new_n933), .A2(new_n934), .A3(new_n677), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT43), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n662), .A2(new_n503), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n650), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n634), .A2(new_n503), .A3(new_n662), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n931), .A2(new_n935), .B1(new_n936), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n936), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n942), .A2(new_n943), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n673), .A2(new_n928), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(KEYINPUT106), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(KEYINPUT106), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  NAND4_X1  g0751(.A1(new_n944), .A2(new_n948), .A3(new_n949), .A4(new_n945), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n928), .A2(new_n678), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(KEYINPUT45), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(KEYINPUT45), .ZN(new_n956));
  AND2_X1   g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n928), .A2(new_n678), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT44), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n928), .A2(KEYINPUT44), .A3(new_n678), .ZN(new_n961));
  AND2_X1   g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n674), .B1(new_n957), .B2(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n955), .A2(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n673), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n675), .A2(new_n661), .A3(new_n663), .ZN(new_n967));
  OR2_X1    g0767(.A1(new_n967), .A2(KEYINPUT108), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n967), .A2(KEYINPUT108), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n968), .A2(new_n929), .A3(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n724), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n722), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n722), .B1(new_n966), .B2(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(KEYINPUT107), .B(KEYINPUT41), .Z(new_n974));
  XOR2_X1   g0774(.A(new_n681), .B(new_n974), .Z(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n727), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n940), .A2(new_n741), .ZN(new_n978));
  INV_X1    g0778(.A(G311), .ZN(new_n979));
  OAI22_X1  g0779(.A1(new_n755), .A2(new_n979), .B1(new_n770), .B2(new_n450), .ZN(new_n980));
  XOR2_X1   g0780(.A(new_n980), .B(KEYINPUT109), .Z(new_n981));
  NAND3_X1  g0781(.A1(new_n824), .A2(KEYINPUT46), .A3(G116), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n322), .B1(new_n772), .B2(new_n822), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(G107), .B2(new_n761), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(KEYINPUT110), .B(KEYINPUT46), .Z(new_n986));
  OAI21_X1  g0786(.A(new_n986), .B1(new_n758), .B2(new_n455), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n988), .A2(KEYINPUT111), .ZN(new_n989));
  AOI22_X1  g0789(.A1(G294), .A2(new_n764), .B1(new_n787), .B2(G317), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(KEYINPUT111), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n767), .A2(G97), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n989), .A2(new_n990), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n755), .A2(new_n829), .B1(new_n766), .B2(new_n252), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(G58), .B2(new_n824), .ZN(new_n995));
  INV_X1    g0795(.A(G150), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n770), .A2(new_n996), .B1(new_n760), .B2(new_n242), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(KEYINPUT112), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n322), .B1(new_n787), .B2(G137), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G159), .A2(new_n764), .B1(new_n773), .B2(G50), .ZN(new_n1000));
  NAND4_X1  g0800(.A1(new_n995), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n997), .A2(KEYINPUT112), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n985), .A2(new_n993), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT47), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n747), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n1004), .B2(new_n1003), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n734), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n744), .B1(new_n218), .B2(new_n303), .C1(new_n236), .C2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n728), .A3(new_n1008), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n953), .A2(new_n977), .B1(new_n978), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(KEYINPUT113), .ZN(G387));
  AOI21_X1  g0811(.A(new_n682), .B1(new_n722), .B2(new_n971), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n722), .B2(new_n971), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n971), .A2(new_n727), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1007), .B1(new_n233), .B2(G45), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n683), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1015), .B1(new_n1016), .B2(new_n731), .ZN(new_n1017));
  AOI21_X1  g0817(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n272), .A2(new_n202), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n683), .B(new_n1018), .C1(new_n1019), .C2(KEYINPUT50), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(KEYINPUT50), .B2(new_n1019), .ZN(new_n1021));
  OAI22_X1  g0821(.A1(new_n1017), .A2(new_n1021), .B1(G107), .B2(new_n218), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n729), .B1(new_n1022), .B2(new_n744), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n758), .A2(new_n252), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(G150), .B2(new_n787), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1025), .A2(new_n248), .A3(new_n992), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n755), .A2(new_n784), .B1(new_n770), .B2(new_n202), .ZN(new_n1027));
  OAI22_X1  g0827(.A1(new_n763), .A2(new_n352), .B1(new_n772), .B2(new_n242), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n760), .A2(new_n303), .ZN(new_n1029));
  NOR4_X1   g0829(.A1(new_n1026), .A2(new_n1027), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(G317), .A2(new_n771), .B1(new_n773), .B2(G303), .ZN(new_n1031));
  XOR2_X1   g0831(.A(KEYINPUT114), .B(G322), .Z(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n1031), .B1(new_n979), .B2(new_n763), .C1(new_n755), .C2(new_n1033), .ZN(new_n1034));
  XOR2_X1   g0834(.A(new_n1034), .B(KEYINPUT115), .Z(new_n1035));
  OR2_X1    g0835(.A1(new_n1035), .A2(KEYINPUT48), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(KEYINPUT48), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n824), .A2(G294), .B1(new_n761), .B2(G283), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT49), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n322), .B1(new_n750), .B2(new_n756), .C1(new_n455), .C2(new_n766), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT116), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1030), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1045));
  OAI221_X1 g0845(.A(new_n1023), .B1(new_n664), .B2(new_n741), .C1(new_n1045), .C2(new_n747), .ZN(new_n1046));
  AND2_X1   g0846(.A1(new_n1014), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1013), .A2(new_n1047), .ZN(G393));
  NAND2_X1  g0848(.A1(new_n966), .A2(KEYINPUT117), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT117), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n963), .A2(new_n965), .A3(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n727), .A3(new_n1051), .ZN(new_n1052));
  OAI221_X1 g0852(.A(new_n744), .B1(new_n461), .B2(new_n218), .C1(new_n240), .C2(new_n1007), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(G317), .A2(new_n778), .B1(new_n771), .B2(G311), .ZN(new_n1054));
  XOR2_X1   g0854(.A(new_n1054), .B(KEYINPUT52), .Z(new_n1055));
  OAI221_X1 g0855(.A(new_n322), .B1(new_n760), .B2(new_n455), .C1(new_n496), .C2(new_n766), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1033), .A2(new_n750), .B1(new_n819), .B2(new_n772), .ZN(new_n1057));
  OAI22_X1  g0857(.A1(new_n822), .A2(new_n758), .B1(new_n763), .B2(new_n450), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n755), .A2(new_n996), .B1(new_n770), .B2(new_n784), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT51), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n761), .A2(G77), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1062), .B(new_n248), .C1(new_n209), .C2(new_n766), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n763), .A2(new_n202), .B1(new_n772), .B2(new_n352), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n758), .A2(new_n242), .B1(new_n750), .B2(new_n829), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1055), .A2(new_n1059), .B1(new_n1061), .B2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n728), .B(new_n1053), .C1(new_n1067), .C2(new_n747), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n928), .B2(new_n742), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  AND2_X1   g0870(.A1(new_n966), .A2(new_n972), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n681), .B1(new_n966), .B2(new_n972), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1052), .B(new_n1070), .C1(new_n1071), .C2(new_n1072), .ZN(G390));
  INV_X1    g0873(.A(new_n909), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n384), .A2(new_n806), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n660), .B(new_n1075), .C1(new_n696), .C2(new_n700), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1074), .B1(new_n1076), .B2(new_n805), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n889), .B1(new_n884), .B2(new_n885), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n810), .A2(new_n805), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n889), .B1(new_n1080), .B2(new_n909), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n1077), .A2(new_n1079), .B1(new_n1081), .B2(new_n888), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n720), .A2(new_n809), .A3(new_n909), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(KEYINPUT118), .B1(new_n1082), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1076), .A2(new_n805), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n909), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1087), .A2(new_n1078), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT118), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n882), .B(new_n887), .C1(new_n895), .C2(new_n889), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1088), .A2(new_n1089), .A3(new_n1090), .A4(new_n1083), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n908), .A2(new_n809), .ZN(new_n1092));
  NOR3_X1   g0892(.A1(new_n1092), .A2(new_n1074), .A3(new_n669), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1082), .A2(new_n1093), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1085), .A2(new_n1091), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n909), .B1(new_n720), .B2(new_n809), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1080), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1074), .B1(new_n1092), .B2(new_n669), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1098), .A2(new_n805), .A3(new_n1076), .A4(new_n1083), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n630), .B(new_n917), .C1(new_n702), .C2(new_n439), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1095), .A2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1101), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1105), .A2(new_n1085), .A3(new_n1091), .A4(new_n1094), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1104), .A2(new_n681), .A3(new_n1106), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1085), .A2(new_n1091), .A3(new_n727), .A4(new_n1094), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n728), .B1(new_n817), .B2(new_n272), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n758), .A2(new_n996), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(new_n1110), .B(KEYINPUT53), .ZN(new_n1111));
  XOR2_X1   g0911(.A(KEYINPUT54), .B(G143), .Z(new_n1112));
  AOI22_X1  g0912(.A1(new_n773), .A2(new_n1112), .B1(new_n767), .B2(G50), .ZN(new_n1113));
  INV_X1    g0913(.A(G128), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1111), .B(new_n1113), .C1(new_n1114), .C2(new_n755), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G132), .A2(new_n771), .B1(new_n764), .B2(G137), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n322), .B1(new_n787), .B2(G125), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1116), .B(new_n1117), .C1(new_n784), .C2(new_n760), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(G283), .A2(new_n778), .B1(new_n773), .B2(G97), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1119), .B1(new_n496), .B2(new_n763), .C1(new_n455), .C2(new_n770), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n248), .B1(new_n824), .B2(G87), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n787), .A2(G294), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1121), .A2(new_n1122), .A3(new_n839), .A4(new_n1062), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n1115), .A2(new_n1118), .B1(new_n1120), .B2(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1109), .B1(new_n1124), .B2(new_n743), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1125), .B1(new_n888), .B2(new_n739), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1108), .A2(new_n1126), .ZN(new_n1127));
  AND2_X1   g0927(.A1(new_n1107), .A2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(G378));
  NAND2_X1  g0929(.A1(new_n300), .A2(new_n333), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n295), .A2(new_n861), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1130), .B(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1133), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1132), .B(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1136), .A2(new_n738), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n728), .B1(new_n817), .B2(G50), .ZN(new_n1138));
  INV_X1    g0938(.A(G41), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n322), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1140), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT119), .Z(new_n1142));
  OAI22_X1  g0942(.A1(new_n339), .A2(new_n766), .B1(new_n772), .B2(new_n303), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1143), .A2(new_n1024), .A3(new_n1140), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n761), .A2(G68), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n778), .A2(G116), .B1(new_n787), .B2(G283), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(G97), .A2(new_n764), .B1(new_n771), .B2(G107), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n1144), .A2(new_n1145), .A3(new_n1146), .A4(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT58), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1142), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI22_X1  g0950(.A1(new_n1112), .A2(new_n824), .B1(new_n771), .B2(G128), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n778), .A2(G125), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1151), .B(new_n1152), .C1(new_n996), .C2(new_n760), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(G132), .A2(new_n764), .B1(new_n773), .B2(G137), .ZN(new_n1154));
  OR2_X1    g0954(.A1(new_n1154), .A2(KEYINPUT120), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(KEYINPUT120), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1153), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT59), .ZN(new_n1158));
  AND2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n273), .B(new_n1139), .C1(new_n766), .C2(new_n784), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1160), .B1(G124), .B2(new_n787), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1150), .B1(new_n1149), .B2(new_n1148), .C1(new_n1159), .C2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1138), .B1(new_n1163), .B2(new_n743), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1137), .A2(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1135), .B1(new_n919), .B2(G330), .ZN(new_n1167));
  AND4_X1   g0967(.A1(G330), .A2(new_n912), .A3(new_n1135), .A4(new_n915), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n900), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n919), .A2(G330), .A3(new_n1135), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n916), .A2(new_n1136), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n900), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1170), .A2(new_n1171), .A3(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1169), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1166), .B1(new_n1174), .B2(new_n727), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1106), .A2(new_n1102), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1176), .A2(KEYINPUT57), .A3(new_n1174), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n681), .ZN(new_n1178));
  AOI22_X1  g0978(.A1(new_n1106), .A2(new_n1102), .B1(new_n1173), .B2(new_n1169), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1179), .A2(KEYINPUT57), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1175), .B1(new_n1178), .B2(new_n1180), .ZN(G375));
  NAND3_X1  g0981(.A1(new_n1097), .A2(new_n1101), .A3(new_n1099), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1103), .A2(new_n976), .A3(new_n1182), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n755), .A2(new_n837), .B1(new_n750), .B2(new_n1114), .ZN(new_n1184));
  AOI211_X1 g0984(.A(new_n322), .B(new_n1184), .C1(G58), .C2(new_n767), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G159), .A2(new_n824), .B1(new_n764), .B2(new_n1112), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G137), .A2(new_n771), .B1(new_n773), .B2(G150), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n761), .A2(G50), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n322), .B1(new_n766), .B2(new_n252), .ZN(new_n1190));
  XNOR2_X1  g0990(.A(new_n1190), .B(KEYINPUT121), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n770), .A2(new_n822), .B1(new_n772), .B2(new_n496), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n755), .A2(new_n819), .B1(new_n763), .B2(new_n455), .ZN(new_n1193));
  OR4_X1    g0993(.A1(new_n1029), .A2(new_n1191), .A3(new_n1192), .A4(new_n1193), .ZN(new_n1194));
  OAI22_X1  g0994(.A1(new_n758), .A2(new_n461), .B1(new_n750), .B2(new_n450), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT122), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1189), .B1(new_n1194), .B2(new_n1196), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n747), .B1(new_n1197), .B2(KEYINPUT123), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1198), .B1(KEYINPUT123), .B2(new_n1197), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1199), .B(new_n728), .C1(G68), .C2(new_n817), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(new_n1074), .B2(new_n738), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n1100), .B2(new_n727), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1183), .A2(new_n1202), .ZN(G381));
  INV_X1    g1003(.A(new_n1175), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n682), .B1(new_n1179), .B2(KEYINPUT57), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1176), .A2(new_n1174), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT57), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1204), .B1(new_n1205), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n1128), .ZN(new_n1210));
  INV_X1    g1010(.A(G390), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1013), .A2(new_n793), .A3(new_n1047), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1211), .A2(new_n848), .A3(new_n1213), .ZN(new_n1214));
  NOR4_X1   g1014(.A1(G387), .A2(new_n1210), .A3(G381), .A4(new_n1214), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(new_n1215), .B(KEYINPUT124), .ZN(G407));
  OAI211_X1 g1016(.A(G407), .B(G213), .C1(G343), .C2(new_n1210), .ZN(G409));
  AOI21_X1  g1017(.A(new_n793), .B1(new_n1013), .B2(new_n1047), .ZN(new_n1218));
  OAI21_X1  g1018(.A(G390), .B1(new_n1213), .B2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT113), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1218), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1220), .B1(new_n1221), .B2(new_n1212), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1010), .B(new_n1219), .C1(G390), .C2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(KEYINPUT113), .B1(new_n1213), .B2(new_n1218), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1225), .A2(new_n1211), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1010), .B1(new_n1226), .B2(new_n1219), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1224), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1205), .A2(new_n1208), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1128), .B1(new_n1229), .B2(new_n1175), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT60), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1182), .A2(new_n1231), .ZN(new_n1232));
  NAND4_X1  g1032(.A1(new_n1097), .A2(new_n1101), .A3(new_n1099), .A4(KEYINPUT60), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1232), .A2(new_n1103), .A3(new_n681), .A4(new_n1233), .ZN(new_n1234));
  AND3_X1   g1034(.A1(new_n1234), .A2(new_n848), .A3(new_n1202), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n848), .B1(new_n1234), .B2(new_n1202), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(G213), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1238), .A2(G343), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1175), .A2(new_n1107), .A3(new_n1127), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n1206), .A2(new_n975), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1240), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  NOR3_X1   g1043(.A1(new_n1230), .A2(new_n1237), .A3(new_n1243), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1228), .B1(new_n1244), .B2(KEYINPUT63), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(G375), .A2(G378), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1237), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1175), .A2(new_n1107), .A3(new_n1127), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1179), .A2(new_n976), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1239), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1246), .A2(KEYINPUT63), .A3(new_n1247), .A4(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1234), .A2(new_n1202), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(G384), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1234), .A2(new_n848), .A3(new_n1202), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1253), .A2(G2897), .A3(new_n1254), .A4(new_n1239), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1239), .A2(G2897), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n1230), .B2(new_n1243), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT61), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1251), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(KEYINPUT125), .B1(new_n1245), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1010), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1222), .A2(G390), .ZN(new_n1264));
  AND2_X1   g1064(.A1(new_n1052), .A2(new_n1070), .ZN(new_n1265));
  OR2_X1    g1065(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1266));
  AOI22_X1  g1066(.A1(new_n1265), .A2(new_n1266), .B1(new_n1221), .B2(new_n1212), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1263), .B1(new_n1264), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n1223), .ZN(new_n1269));
  OAI211_X1 g1069(.A(new_n1250), .B(new_n1247), .C1(new_n1128), .C2(new_n1209), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT63), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT125), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1128), .A2(new_n1175), .A3(new_n1249), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1274), .B(new_n1240), .C1(new_n1209), .C2(new_n1128), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT61), .B1(new_n1275), .B2(new_n1258), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1272), .A2(new_n1273), .A3(new_n1276), .A4(new_n1251), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1262), .A2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1270), .A2(KEYINPUT62), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT62), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1246), .A2(new_n1280), .A3(new_n1247), .A4(new_n1250), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1279), .B(new_n1281), .C1(new_n1276), .C2(KEYINPUT126), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1259), .A2(KEYINPUT126), .A3(new_n1260), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1269), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1278), .A2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT127), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1278), .A2(new_n1284), .A3(KEYINPUT127), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(G405));
  NAND2_X1  g1089(.A1(new_n1246), .A2(new_n1210), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(new_n1247), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(new_n1228), .ZN(G402));
endmodule


