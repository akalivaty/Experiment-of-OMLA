//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 0 1 0 0 1 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:44 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  INV_X1    g000(.A(KEYINPUT69), .ZN(new_n187));
  XOR2_X1   g001(.A(KEYINPUT68), .B(KEYINPUT32), .Z(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  NOR2_X1   g003(.A1(G237), .A2(G953), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G210), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n191), .B(KEYINPUT27), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT26), .B(G101), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G143), .ZN(new_n199));
  AOI211_X1 g013(.A(new_n196), .B(new_n198), .C1(new_n199), .C2(G146), .ZN(new_n200));
  INV_X1    g014(.A(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(G128), .B1(new_n196), .B2(new_n197), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n195), .A2(KEYINPUT64), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT64), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  AOI21_X1  g020(.A(G146), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(G143), .ZN(new_n209));
  OAI211_X1 g023(.A(new_n202), .B(new_n203), .C1(new_n207), .C2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n209), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n212), .B1(new_n199), .B2(G146), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n203), .B1(new_n213), .B2(new_n202), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n201), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  INV_X1    g030(.A(G134), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(G137), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI211_X1 g034(.A(KEYINPUT65), .B(new_n216), .C1(new_n217), .C2(G137), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G131), .ZN(new_n223));
  INV_X1    g037(.A(G137), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(KEYINPUT11), .A3(G134), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n217), .A2(G137), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n222), .A2(new_n223), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n224), .A2(G134), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n226), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G131), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n221), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT65), .B1(new_n230), .B2(new_n216), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n228), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G131), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n229), .ZN(new_n239));
  AND2_X1   g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n196), .B1(new_n199), .B2(G146), .ZN(new_n243));
  AOI22_X1  g057(.A1(new_n213), .A2(new_n242), .B1(new_n243), .B2(new_n240), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n215), .A2(new_n234), .B1(new_n239), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G116), .B(G119), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(KEYINPUT2), .B(G113), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g063(.A(KEYINPUT2), .B(G113), .Z(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(new_n246), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n245), .A2(new_n253), .ZN(new_n254));
  AOI211_X1 g068(.A(G131), .B(new_n227), .C1(new_n220), .C2(new_n221), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n223), .B1(new_n222), .B2(new_n228), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n244), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n207), .A2(new_n209), .ZN(new_n258));
  INV_X1    g072(.A(new_n202), .ZN(new_n259));
  OAI21_X1  g073(.A(KEYINPUT66), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n200), .B1(new_n260), .B2(new_n210), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n257), .B1(new_n261), .B2(new_n233), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(new_n252), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT28), .B1(new_n254), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n215), .A2(new_n234), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n265), .A2(new_n253), .A3(new_n257), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT28), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n194), .B1(new_n264), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT31), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n252), .B1(new_n245), .B2(KEYINPUT30), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n257), .B(KEYINPUT30), .C1(new_n261), .C2(new_n233), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT67), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n265), .A2(KEYINPUT67), .A3(KEYINPUT30), .A4(new_n257), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n271), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n266), .A2(new_n194), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n270), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n274), .A2(new_n275), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT30), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n253), .B1(new_n262), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n277), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n282), .A2(KEYINPUT31), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n269), .B1(new_n278), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(G472), .A2(G902), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n187), .B(new_n189), .C1(new_n285), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n264), .A2(new_n268), .ZN(new_n289));
  INV_X1    g103(.A(new_n194), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n194), .B1(new_n282), .B2(new_n266), .ZN(new_n292));
  NOR3_X1   g106(.A1(new_n291), .A2(new_n292), .A3(KEYINPUT29), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  OR2_X1    g108(.A1(new_n268), .A2(KEYINPUT70), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n268), .A2(KEYINPUT70), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n264), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n194), .A2(KEYINPUT29), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  OAI21_X1  g113(.A(G472), .B1(new_n293), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n278), .A2(new_n284), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n289), .A2(new_n290), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n287), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(KEYINPUT69), .B1(new_n303), .B2(KEYINPUT32), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n303), .A2(new_n188), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n288), .B(new_n300), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(G214), .B1(G237), .B2(G902), .ZN(new_n307));
  OAI21_X1  g121(.A(G210), .B1(G237), .B2(G902), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT82), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  XNOR2_X1  g124(.A(G110), .B(G122), .ZN(new_n311));
  INV_X1    g125(.A(G104), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT3), .B1(new_n312), .B2(G107), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT3), .ZN(new_n314));
  INV_X1    g128(.A(G107), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n314), .A2(new_n315), .A3(G104), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n312), .A2(G107), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G101), .ZN(new_n319));
  INV_X1    g133(.A(G101), .ZN(new_n320));
  NAND4_X1  g134(.A1(new_n313), .A2(new_n316), .A3(new_n320), .A4(new_n317), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(KEYINPUT4), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT4), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n318), .A2(new_n323), .A3(G101), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n252), .A3(new_n324), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n325), .A2(KEYINPUT79), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n322), .A2(new_n252), .A3(new_n327), .A4(new_n324), .ZN(new_n328));
  INV_X1    g142(.A(new_n317), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n312), .A2(G107), .ZN(new_n330));
  OAI21_X1  g144(.A(G101), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n321), .ZN(new_n332));
  INV_X1    g146(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n246), .A2(KEYINPUT5), .ZN(new_n334));
  INV_X1    g148(.A(G116), .ZN(new_n335));
  OR3_X1    g149(.A1(new_n335), .A2(KEYINPUT5), .A3(G119), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(G113), .A3(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(new_n251), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n328), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT80), .B1(new_n326), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n325), .A2(KEYINPUT79), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT80), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n341), .A2(new_n342), .A3(new_n328), .A4(new_n338), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n311), .B1(new_n340), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n311), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n326), .A2(new_n339), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT6), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n339), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n342), .B1(new_n348), .B2(new_n341), .ZN(new_n349));
  INV_X1    g163(.A(new_n343), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n345), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT6), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n347), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n244), .A2(G125), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n261), .B2(G125), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G224), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(G953), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n359), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n354), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT7), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n357), .B1(new_n365), .B2(new_n359), .ZN(new_n366));
  INV_X1    g180(.A(new_n346), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n356), .A2(KEYINPUT7), .A3(new_n361), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n337), .A2(new_n251), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n332), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n338), .ZN(new_n371));
  XOR2_X1   g185(.A(KEYINPUT81), .B(KEYINPUT8), .Z(new_n372));
  XNOR2_X1  g186(.A(new_n372), .B(new_n311), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n366), .A2(new_n367), .A3(new_n368), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n294), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n310), .B1(new_n364), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n363), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n379), .B1(new_n347), .B2(new_n353), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n380), .A2(new_n309), .A3(new_n376), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n307), .B1(new_n378), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(G110), .B(G140), .ZN(new_n383));
  INV_X1    g197(.A(G953), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G227), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n383), .B(new_n385), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT1), .B1(new_n199), .B2(G146), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n243), .B1(G128), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n333), .B1(new_n388), .B2(new_n200), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT10), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n332), .A2(new_n390), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n215), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n244), .A2(new_n324), .A3(new_n322), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n391), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n255), .A2(new_n256), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(KEYINPUT77), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT77), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n239), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n386), .B1(new_n395), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n395), .A2(new_n239), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n395), .A2(new_n400), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT12), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n201), .B(new_n332), .C1(new_n211), .C2(new_n214), .ZN(new_n407));
  AOI211_X1 g221(.A(new_n406), .B(new_n396), .C1(new_n407), .C2(new_n389), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n389), .ZN(new_n409));
  AOI21_X1  g223(.A(KEYINPUT12), .B1(new_n409), .B2(new_n239), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT78), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n408), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n396), .B1(new_n407), .B2(new_n389), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT78), .B1(new_n413), .B2(KEYINPUT12), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n405), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(G469), .B(new_n404), .C1(new_n415), .C2(new_n386), .ZN(new_n416));
  INV_X1    g230(.A(G469), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n401), .B1(new_n412), .B2(new_n414), .ZN(new_n418));
  AOI22_X1  g232(.A1(new_n390), .A2(new_n389), .B1(new_n215), .B2(new_n392), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n419), .A2(new_n394), .A3(new_n399), .A4(new_n397), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n386), .B1(new_n420), .B2(new_n403), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n417), .B(new_n294), .C1(new_n418), .C2(new_n421), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n417), .A2(new_n294), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n416), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n384), .A2(G952), .ZN(new_n426));
  NAND2_X1  g240(.A1(G234), .A2(G237), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(G902), .A3(G953), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(G898), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n429), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT92), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n199), .A2(G128), .ZN(new_n435));
  INV_X1    g249(.A(G128), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(G143), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G134), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n435), .A2(new_n217), .A3(new_n437), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(G122), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n442), .A2(G116), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT14), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n442), .A2(G116), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n443), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n446), .B1(new_n444), .B2(new_n443), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n335), .A2(G122), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT89), .B1(new_n448), .B2(new_n443), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n335), .A2(G122), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT89), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n445), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(G107), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n453), .A2(KEYINPUT91), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(KEYINPUT91), .ZN(new_n455));
  OAI221_X1 g269(.A(new_n441), .B1(new_n315), .B2(new_n447), .C1(new_n454), .C2(new_n455), .ZN(new_n456));
  AND3_X1   g270(.A1(new_n449), .A2(G107), .A3(new_n452), .ZN(new_n457));
  XOR2_X1   g271(.A(KEYINPUT90), .B(KEYINPUT13), .Z(new_n458));
  AND3_X1   g272(.A1(new_n435), .A2(new_n437), .A3(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(G134), .B1(new_n435), .B2(new_n458), .ZN(new_n460));
  OAI221_X1 g274(.A(new_n440), .B1(new_n457), .B2(new_n453), .C1(new_n459), .C2(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT9), .B(G234), .ZN(new_n462));
  INV_X1    g276(.A(G217), .ZN(new_n463));
  NOR3_X1   g277(.A1(new_n462), .A2(new_n463), .A3(G953), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n456), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n464), .B1(new_n456), .B2(new_n461), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n434), .B1(new_n467), .B2(G902), .ZN(new_n468));
  INV_X1    g282(.A(G478), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(KEYINPUT15), .ZN(new_n470));
  INV_X1    g284(.A(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n456), .A2(new_n461), .ZN(new_n472));
  INV_X1    g286(.A(new_n464), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n456), .A2(new_n461), .A3(new_n464), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n476), .A2(KEYINPUT92), .A3(new_n294), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n468), .A2(new_n471), .A3(new_n477), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n476), .A2(KEYINPUT92), .A3(new_n294), .A4(new_n470), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n433), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  XOR2_X1   g294(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(G113), .B(G122), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(new_n312), .ZN(new_n484));
  INV_X1    g298(.A(G140), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G125), .ZN(new_n486));
  INV_X1    g300(.A(G125), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(G140), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT87), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n489), .A2(new_n490), .A3(KEYINPUT19), .ZN(new_n491));
  XOR2_X1   g305(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n492));
  OAI21_X1  g306(.A(new_n491), .B1(new_n489), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n208), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT16), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n485), .A3(G125), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT73), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n496), .B(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT72), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n489), .A2(new_n499), .A3(KEYINPUT16), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n486), .A2(new_n488), .ZN(new_n501));
  OAI21_X1  g315(.A(KEYINPUT72), .B1(new_n501), .B2(new_n495), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n498), .A2(new_n500), .A3(G146), .A4(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n494), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n190), .A2(G143), .A3(G214), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT86), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n505), .B(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(G237), .ZN(new_n508));
  AND4_X1   g322(.A1(KEYINPUT84), .A2(new_n508), .A3(new_n384), .A4(G214), .ZN(new_n509));
  AOI21_X1  g323(.A(KEYINPUT84), .B1(new_n190), .B2(G214), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n199), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT85), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT85), .B(new_n199), .C1(new_n509), .C2(new_n510), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n507), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n515), .A2(new_n223), .ZN(new_n516));
  AOI211_X1 g330(.A(G131), .B(new_n507), .C1(new_n513), .C2(new_n514), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n504), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n507), .ZN(new_n519));
  INV_X1    g333(.A(new_n514), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n508), .A2(new_n384), .A3(G214), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT84), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n190), .A2(KEYINPUT84), .A3(G214), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g339(.A(KEYINPUT85), .B1(new_n525), .B2(new_n199), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n519), .B1(new_n520), .B2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n527), .A2(KEYINPUT18), .A3(G131), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n501), .B(new_n208), .ZN(new_n529));
  NAND2_X1  g343(.A1(KEYINPUT18), .A2(G131), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n529), .B1(new_n515), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n484), .B1(new_n518), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n498), .A2(new_n500), .A3(new_n502), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(new_n208), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n503), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n536), .B1(new_n516), .B2(KEYINPUT17), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n527), .A2(G131), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT17), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n515), .A2(new_n223), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n537), .A2(new_n541), .B1(new_n528), .B2(new_n531), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n533), .B1(new_n484), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g357(.A1(G475), .A2(G902), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n544), .B(KEYINPUT88), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n482), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NOR3_X1   g360(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT17), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n535), .A2(new_n503), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n538), .B2(new_n539), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n484), .B(new_n532), .C1(new_n547), .C2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n484), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n528), .A2(new_n531), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n494), .A2(new_n503), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n538), .B2(new_n540), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n551), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT20), .ZN(new_n557));
  INV_X1    g371(.A(new_n545), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n550), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n537), .A2(new_n541), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n484), .B1(new_n561), .B2(new_n532), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n294), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n546), .A2(new_n559), .B1(new_n563), .B2(G475), .ZN(new_n564));
  OAI21_X1  g378(.A(G221), .B1(new_n462), .B2(G902), .ZN(new_n565));
  NAND4_X1  g379(.A1(new_n425), .A2(new_n480), .A3(new_n564), .A4(new_n565), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n382), .A2(new_n566), .ZN(new_n567));
  OAI211_X1 g381(.A(KEYINPUT71), .B(KEYINPUT23), .C1(new_n436), .C2(G119), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n436), .B(G119), .C1(KEYINPUT71), .C2(KEYINPUT23), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G110), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT24), .B(G110), .Z(new_n572));
  XNOR2_X1  g386(.A(G119), .B(G128), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n575), .B1(new_n535), .B2(new_n503), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n489), .A2(new_n208), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n570), .A2(G110), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n572), .A2(new_n573), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n503), .B(new_n577), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g395(.A(KEYINPUT74), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n536), .A2(new_n574), .A3(new_n571), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT74), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n584), .A3(new_n580), .ZN(new_n585));
  XOR2_X1   g399(.A(KEYINPUT22), .B(G137), .Z(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(KEYINPUT75), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n384), .A2(G221), .A3(G234), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n587), .B(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n582), .A2(new_n585), .A3(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n583), .A2(new_n580), .A3(new_n589), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n463), .B1(G234), .B2(new_n294), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(G902), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n595), .B(KEYINPUT76), .Z(new_n596));
  NOR2_X1   g410(.A1(new_n593), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT25), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n591), .A2(new_n592), .A3(new_n598), .A4(new_n294), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n594), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n591), .A2(new_n592), .A3(new_n294), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(KEYINPUT25), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n597), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n306), .A2(new_n567), .A3(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(G101), .ZN(G3));
  INV_X1    g420(.A(new_n307), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n364), .A2(new_n310), .A3(new_n377), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n309), .B1(new_n380), .B2(new_n376), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n433), .ZN(new_n611));
  NOR3_X1   g425(.A1(new_n467), .A2(G478), .A3(G902), .ZN(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(KEYINPUT33), .B1(new_n465), .B2(new_n466), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n474), .A2(new_n615), .A3(new_n475), .ZN(new_n616));
  AOI21_X1  g430(.A(G902), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n613), .B1(new_n617), .B2(new_n469), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n564), .A2(new_n618), .ZN(new_n619));
  AND3_X1   g433(.A1(new_n610), .A2(new_n611), .A3(new_n619), .ZN(new_n620));
  AND2_X1   g434(.A1(new_n425), .A2(new_n565), .ZN(new_n621));
  NAND2_X1  g435(.A1(KEYINPUT93), .A2(G472), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n285), .B2(G902), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT31), .B1(new_n282), .B2(new_n283), .ZN(new_n625));
  AOI211_X1 g439(.A(new_n270), .B(new_n277), .C1(new_n279), .C2(new_n281), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n302), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(new_n294), .A3(new_n622), .ZN(new_n628));
  AND3_X1   g442(.A1(new_n624), .A2(new_n628), .A3(new_n604), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n620), .A2(new_n621), .A3(new_n629), .ZN(new_n630));
  XOR2_X1   g444(.A(new_n630), .B(KEYINPUT94), .Z(new_n631));
  XNOR2_X1  g445(.A(KEYINPUT34), .B(G104), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  XOR2_X1   g447(.A(new_n433), .B(KEYINPUT96), .Z(new_n634));
  NAND2_X1  g448(.A1(new_n610), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT95), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n481), .B1(new_n556), .B2(new_n558), .ZN(new_n637));
  AOI211_X1 g451(.A(new_n545), .B(new_n482), .C1(new_n550), .C2(new_n555), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n556), .A2(new_n558), .A3(new_n481), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n546), .A2(KEYINPUT95), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n563), .A2(G475), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n478), .A2(new_n479), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n642), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n635), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(new_n621), .A3(new_n629), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  AND2_X1   g464(.A1(new_n582), .A2(new_n585), .ZN(new_n651));
  OR2_X1    g465(.A1(new_n590), .A2(KEYINPUT36), .ZN(new_n652));
  OR2_X1    g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n651), .A2(new_n652), .ZN(new_n654));
  INV_X1    g468(.A(new_n596), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n653), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n603), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n656), .B1(new_n657), .B2(new_n600), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n624), .A2(new_n628), .A3(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT97), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n624), .A2(new_n628), .A3(new_n658), .A4(KEYINPUT97), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n567), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT37), .B(G110), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G12));
  OAI21_X1  g480(.A(new_n428), .B1(G900), .B2(new_n430), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n642), .A2(new_n643), .A3(new_n645), .A4(new_n667), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n307), .B(new_n658), .C1(new_n378), .C2(new_n381), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n306), .A3(new_n621), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT98), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n670), .A2(new_n306), .A3(KEYINPUT98), .A4(new_n621), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  XNOR2_X1  g490(.A(new_n667), .B(KEYINPUT39), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n621), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(new_n678), .B(KEYINPUT40), .Z(new_n679));
  NAND2_X1  g493(.A1(new_n608), .A2(new_n609), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT38), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n276), .A2(new_n277), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n254), .A2(new_n263), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n682), .B1(new_n290), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g498(.A(G472), .B1(new_n684), .B2(G902), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n288), .B(new_n685), .C1(new_n304), .C2(new_n305), .ZN(new_n686));
  NOR4_X1   g500(.A1(new_n658), .A2(new_n564), .A3(new_n644), .A4(new_n607), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n679), .A2(new_n681), .A3(new_n686), .A4(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n688), .B(new_n199), .Z(G45));
  AND3_X1   g503(.A1(new_n610), .A2(new_n619), .A3(new_n667), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n690), .A2(new_n306), .A3(new_n621), .A4(new_n658), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G146), .ZN(G48));
  NAND2_X1  g506(.A1(new_n410), .A2(new_n411), .ZN(new_n693));
  INV_X1    g507(.A(new_n408), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n693), .A2(new_n414), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n420), .A2(new_n403), .ZN(new_n696));
  INV_X1    g510(.A(new_n386), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n695), .A2(new_n402), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(G469), .B1(new_n698), .B2(G902), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n565), .A3(new_n422), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT99), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n699), .A2(KEYINPUT99), .A3(new_n565), .A4(new_n422), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n620), .A2(new_n306), .A3(new_n704), .A4(new_n604), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT100), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G15));
  NAND4_X1  g522(.A1(new_n647), .A2(new_n604), .A3(new_n306), .A4(new_n704), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G116), .ZN(G18));
  AND3_X1   g524(.A1(new_n610), .A2(new_n702), .A3(new_n703), .ZN(new_n711));
  AND3_X1   g525(.A1(new_n658), .A2(new_n564), .A3(new_n480), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n306), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  AND3_X1   g528(.A1(new_n680), .A2(new_n307), .A3(new_n634), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n564), .A2(new_n644), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n297), .A2(new_n290), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n301), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n286), .ZN(new_n719));
  OAI21_X1  g533(.A(G472), .B1(new_n285), .B2(G902), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n719), .A2(new_n720), .A3(new_n604), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n704), .A2(new_n715), .A3(new_n716), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  NAND2_X1  g537(.A1(new_n619), .A2(new_n667), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n719), .A2(new_n720), .A3(new_n658), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n711), .A2(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT101), .B(G125), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G27));
  INV_X1    g543(.A(KEYINPUT32), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n730), .B1(new_n285), .B2(new_n287), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n627), .A2(KEYINPUT32), .A3(new_n286), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n731), .A2(new_n732), .A3(KEYINPUT103), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n300), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT103), .B1(new_n731), .B2(new_n732), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n604), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT102), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n422), .B(new_n424), .C1(new_n416), .C2(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n401), .B1(new_n239), .B2(new_n395), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n695), .A2(new_n420), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n739), .B1(new_n740), .B2(new_n697), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT102), .B1(new_n741), .B2(G469), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n565), .B1(new_n738), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n608), .A2(new_n307), .A3(new_n609), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n724), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT42), .B1(new_n736), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n724), .A2(KEYINPUT42), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(new_n306), .A3(new_n745), .A4(new_n604), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n223), .ZN(G33));
  INV_X1    g566(.A(new_n668), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n306), .A2(new_n745), .A3(new_n604), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n741), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n404), .B1(new_n415), .B2(new_n386), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT45), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(G469), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(KEYINPUT46), .A3(new_n424), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n422), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT104), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n762), .A2(KEYINPUT104), .A3(new_n422), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT46), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n767), .B(G469), .C1(new_n760), .C2(G902), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n769), .A2(new_n565), .A3(new_n677), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT105), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n617), .A2(new_n469), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n612), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n564), .ZN(new_n774));
  XOR2_X1   g588(.A(new_n774), .B(KEYINPUT43), .Z(new_n775));
  NAND2_X1  g589(.A1(new_n624), .A2(new_n628), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n776), .A2(new_n658), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n775), .A2(KEYINPUT44), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n744), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT44), .B1(new_n775), .B2(new_n777), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT105), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n769), .A2(new_n783), .A3(new_n565), .A4(new_n677), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n771), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT106), .B(G137), .Z(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(G39));
  NOR4_X1   g601(.A1(new_n306), .A2(new_n604), .A3(new_n724), .A4(new_n744), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(KEYINPUT107), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n769), .A2(KEYINPUT47), .A3(new_n565), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT47), .B1(new_n769), .B2(new_n565), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n789), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT108), .ZN(new_n793));
  INV_X1    g607(.A(KEYINPUT108), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n794), .B(new_n789), .C1(new_n790), .C2(new_n791), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  AND3_X1   g611(.A1(new_n705), .A2(new_n722), .A3(new_n713), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n715), .A2(new_n621), .A3(new_n619), .A4(new_n629), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n605), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(KEYINPUT110), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n605), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n798), .A2(new_n801), .A3(new_n709), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n726), .A2(new_n745), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n754), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n642), .A2(new_n643), .A3(new_n644), .A4(new_n667), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n807), .A2(new_n744), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n808), .A2(new_n306), .A3(new_n621), .A4(new_n658), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n806), .A2(new_n748), .A3(new_n750), .A4(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n564), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n811), .A2(new_n644), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n715), .A2(new_n621), .A3(new_n629), .A4(new_n812), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n664), .A2(KEYINPUT111), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(KEYINPUT111), .B1(new_n664), .B2(new_n813), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n804), .A2(new_n810), .A3(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n691), .A2(new_n727), .ZN(new_n818));
  INV_X1    g632(.A(new_n667), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n743), .A2(new_n658), .A3(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n820), .A2(new_n610), .A3(new_n686), .A4(new_n716), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n675), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT113), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT52), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n822), .A2(new_n823), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n824), .B1(new_n822), .B2(new_n823), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n817), .B(KEYINPUT53), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n822), .A2(KEYINPUT52), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n675), .A2(new_n818), .A3(new_n824), .A4(new_n821), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n809), .A2(new_n754), .A3(new_n805), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n751), .A2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(new_n815), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n664), .A2(KEYINPUT111), .A3(new_n813), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n705), .A2(new_n709), .A3(new_n713), .A4(new_n722), .ZN(new_n837));
  INV_X1    g651(.A(new_n803), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n802), .B1(new_n605), .B2(new_n799), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n833), .A2(new_n836), .A3(new_n837), .A4(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n828), .B1(new_n831), .B2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n827), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n831), .A2(new_n841), .A3(new_n828), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n817), .B(KEYINPUT112), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n826), .B2(new_n825), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n845), .B1(new_n847), .B2(new_n828), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n844), .B1(new_n848), .B2(new_n843), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n774), .B(KEYINPUT43), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n428), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n851), .A2(new_n721), .ZN(new_n852));
  OR2_X1    g666(.A1(new_n790), .A2(new_n791), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n699), .A2(new_n422), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n854), .A2(new_n565), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n779), .B(new_n852), .C1(new_n853), .C2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n681), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n852), .A2(new_n607), .A3(new_n857), .A4(new_n704), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT50), .Z(new_n859));
  AND2_X1   g673(.A1(new_n704), .A2(new_n779), .ZN(new_n860));
  INV_X1    g674(.A(new_n686), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n860), .A2(new_n604), .A3(new_n429), .A4(new_n861), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n862), .A2(new_n811), .A3(new_n773), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n851), .A2(new_n860), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n725), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n856), .A2(new_n859), .A3(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n864), .A2(new_n736), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT48), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n852), .A2(new_n711), .ZN(new_n872));
  INV_X1    g686(.A(new_n619), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n872), .B(new_n426), .C1(new_n873), .C2(new_n862), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n875), .B1(new_n867), .B2(new_n868), .ZN(new_n876));
  OR2_X1    g690(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n849), .A2(new_n877), .B1(G952), .B2(G953), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n854), .B(KEYINPUT49), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n604), .A2(new_n307), .A3(new_n565), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n879), .A2(new_n774), .A3(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n881), .A2(new_n857), .A3(new_n861), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT109), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n878), .A2(new_n883), .ZN(G75));
  AOI21_X1  g698(.A(new_n294), .B1(new_n827), .B2(new_n842), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n309), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n354), .B(KEYINPUT114), .ZN(new_n889));
  INV_X1    g703(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n886), .A2(new_n887), .A3(new_n889), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n363), .B(KEYINPUT55), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n893), .B1(new_n891), .B2(new_n892), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n384), .A2(G952), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n896), .B(KEYINPUT115), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n894), .A2(new_n895), .A3(new_n898), .ZN(G51));
  AOI211_X1 g713(.A(new_n294), .B(new_n761), .C1(new_n827), .C2(new_n842), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n843), .B1(new_n827), .B2(new_n842), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n844), .B1(new_n901), .B2(KEYINPUT116), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT116), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n827), .A2(new_n842), .A3(new_n903), .A4(new_n843), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n423), .B(KEYINPUT57), .Z(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n698), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n900), .B1(new_n908), .B2(KEYINPUT117), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT117), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n906), .B1(new_n902), .B2(new_n904), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n910), .B1(new_n911), .B2(new_n698), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n896), .B1(new_n909), .B2(new_n912), .ZN(G54));
  NAND3_X1  g727(.A1(new_n885), .A2(KEYINPUT58), .A3(G475), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n896), .B1(new_n914), .B2(new_n543), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n543), .B2(new_n914), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT118), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(G60));
  NAND2_X1  g732(.A1(new_n614), .A2(new_n616), .ZN(new_n919));
  NAND2_X1  g733(.A1(G478), .A2(G902), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT59), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n919), .B1(new_n849), .B2(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n905), .A2(new_n919), .A3(new_n921), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n922), .A2(new_n898), .A3(new_n923), .ZN(G63));
  INV_X1    g738(.A(KEYINPUT61), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n925), .A2(KEYINPUT119), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n827), .A2(new_n842), .ZN(new_n927));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT60), .Z(new_n929));
  NAND2_X1  g743(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n898), .B1(new_n930), .B2(new_n593), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n927), .A2(new_n653), .A3(new_n654), .A4(new_n929), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n926), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n925), .A2(KEYINPUT119), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n933), .B(new_n934), .Z(G66));
  NOR3_X1   g749(.A1(new_n432), .A2(new_n358), .A3(new_n384), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n804), .A2(new_n816), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n936), .B1(new_n937), .B2(new_n384), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n890), .B1(G898), .B2(new_n384), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G69));
  OAI21_X1  g754(.A(new_n279), .B1(KEYINPUT30), .B2(new_n245), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(new_n493), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n942), .B(KEYINPUT120), .Z(new_n943));
  AND2_X1   g757(.A1(new_n675), .A2(new_n818), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n688), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT62), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n945), .B(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n812), .A2(new_n619), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n948), .A2(new_n678), .A3(new_n744), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n949), .A2(new_n604), .A3(new_n306), .ZN(new_n950));
  AOI21_X1  g764(.A(KEYINPUT121), .B1(new_n785), .B2(new_n950), .ZN(new_n951));
  AND3_X1   g765(.A1(new_n785), .A2(KEYINPUT121), .A3(new_n950), .ZN(new_n952));
  OAI211_X1 g766(.A(new_n947), .B(new_n796), .C1(new_n951), .C2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n943), .B1(new_n953), .B2(new_n384), .ZN(new_n954));
  OR4_X1    g768(.A1(new_n382), .A2(new_n736), .A3(new_n564), .A4(new_n644), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n771), .A2(new_n784), .A3(new_n956), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n748), .A2(new_n750), .A3(new_n754), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n961));
  AND3_X1   g775(.A1(new_n785), .A2(new_n961), .A3(new_n944), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n961), .B1(new_n785), .B2(new_n944), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n796), .B(new_n960), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT123), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n785), .A2(new_n944), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT122), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n785), .A2(new_n961), .A3(new_n944), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT123), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n959), .B1(new_n795), .B2(new_n793), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n965), .A2(new_n384), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n942), .B1(G900), .B2(G953), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n954), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n384), .B1(G227), .B2(G900), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n975), .A2(KEYINPUT124), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(KEYINPUT124), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n976), .A2(KEYINPUT124), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n977), .A2(new_n980), .ZN(G72));
  NAND2_X1  g795(.A1(G472), .A2(G902), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n982), .B(KEYINPUT126), .ZN(new_n983));
  XNOR2_X1  g797(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT127), .Z(new_n986));
  INV_X1    g800(.A(new_n937), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n986), .B1(new_n953), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n282), .A2(new_n266), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n988), .A2(new_n989), .A3(new_n194), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n985), .B1(new_n292), .B2(new_n682), .ZN(new_n991));
  OAI221_X1 g805(.A(new_n990), .B1(G952), .B2(new_n384), .C1(new_n848), .C2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n965), .A2(new_n937), .A3(new_n972), .ZN(new_n993));
  AOI211_X1 g807(.A(new_n989), .B(new_n194), .C1(new_n993), .C2(new_n986), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n992), .A2(new_n994), .ZN(G57));
endmodule


