//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 0 1 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:43 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n787, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n982, new_n983, new_n984;
  INV_X1    g000(.A(KEYINPUT88), .ZN(new_n202));
  INV_X1    g001(.A(G183gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT27), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT27), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT28), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT27), .B(G183gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n211), .A2(KEYINPUT28), .A3(new_n207), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT66), .ZN(new_n214));
  INV_X1    g013(.A(G169gat), .ZN(new_n215));
  INV_X1    g014(.A(G176gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n214), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT26), .ZN(new_n218));
  OAI21_X1  g017(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n220), .A2(new_n223), .B1(G183gat), .B2(G190gat), .ZN(new_n224));
  AND2_X1   g023(.A1(new_n213), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(G176gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n228), .A2(new_n215), .ZN(new_n229));
  NAND2_X1  g028(.A1(KEYINPUT64), .A2(G169gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n227), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n232));
  NAND2_X1  g031(.A1(G183gat), .A2(G190gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(KEYINPUT24), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(G183gat), .A3(G190gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n203), .A2(new_n207), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n222), .A2(KEYINPUT23), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n215), .A2(new_n216), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT65), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n227), .A2(new_n229), .A3(new_n243), .A4(new_n230), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n232), .A2(new_n239), .A3(new_n242), .A4(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT25), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n217), .A2(KEYINPUT23), .A3(new_n219), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n246), .B1(new_n240), .B2(new_n241), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n203), .A2(KEYINPUT24), .ZN(new_n249));
  AOI22_X1  g048(.A1(new_n249), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n233), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n203), .A2(new_n207), .A3(KEYINPUT67), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT67), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n252), .B1(G183gat), .B2(G190gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n247), .B(new_n248), .C1(new_n250), .C2(new_n254), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n245), .A2(new_n246), .B1(new_n255), .B2(KEYINPUT68), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n237), .A2(new_n253), .A3(new_n251), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT68), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n257), .A2(new_n258), .A3(new_n247), .A4(new_n248), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n225), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G226gat), .A2(G233gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  XOR2_X1   g061(.A(KEYINPUT74), .B(KEYINPUT29), .Z(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NOR3_X1   g063(.A1(new_n260), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT75), .ZN(new_n266));
  AOI211_X1 g065(.A(new_n266), .B(new_n225), .C1(new_n256), .C2(new_n259), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n245), .A2(new_n246), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n255), .A2(KEYINPUT68), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n268), .A2(new_n259), .A3(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n225), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT75), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n267), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n265), .B1(new_n273), .B2(new_n262), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n275));
  OR2_X1    g074(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n275), .A2(KEYINPUT73), .ZN(new_n277));
  XNOR2_X1  g076(.A(G197gat), .B(G204gat), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G211gat), .B(G218gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n274), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G8gat), .B(G36gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(G64gat), .B(G92gat), .ZN(new_n284));
  XOR2_X1   g083(.A(new_n283), .B(new_n284), .Z(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT30), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT77), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT76), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n270), .A2(new_n271), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(new_n266), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n260), .A2(KEYINPUT75), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT29), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n289), .B1(new_n293), .B2(new_n262), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n295), .B1(new_n267), .B2(new_n272), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(KEYINPUT76), .A3(new_n261), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n290), .A2(new_n262), .ZN(new_n299));
  INV_X1    g098(.A(new_n281), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n288), .B1(new_n298), .B2(new_n302), .ZN(new_n303));
  AOI211_X1 g102(.A(KEYINPUT77), .B(new_n301), .C1(new_n294), .C2(new_n297), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n282), .B(new_n287), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n282), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n296), .A2(KEYINPUT76), .A3(new_n261), .ZN(new_n307));
  AOI21_X1  g106(.A(KEYINPUT76), .B1(new_n296), .B2(new_n261), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n302), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT77), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n298), .A2(new_n288), .A3(new_n302), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n306), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n305), .B1(new_n312), .B2(new_n285), .ZN(new_n313));
  XNOR2_X1  g112(.A(KEYINPUT78), .B(KEYINPUT30), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n314), .B1(new_n312), .B2(new_n285), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n202), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n282), .B(new_n285), .C1(new_n303), .C2(new_n304), .ZN(new_n317));
  INV_X1    g116(.A(new_n314), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n282), .B1(new_n303), .B2(new_n304), .ZN(new_n320));
  INV_X1    g119(.A(new_n285), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n319), .A2(new_n322), .A3(KEYINPUT88), .A4(new_n305), .ZN(new_n323));
  XOR2_X1   g122(.A(G1gat), .B(G29gat), .Z(new_n324));
  XNOR2_X1  g123(.A(G57gat), .B(G85gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT83), .B(KEYINPUT0), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT71), .ZN(new_n329));
  XNOR2_X1  g128(.A(G127gat), .B(G134gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT1), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT70), .ZN(new_n332));
  INV_X1    g131(.A(G120gat), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n333), .A3(G113gat), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n330), .A2(new_n331), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G113gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(G120gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n333), .A2(G113gat), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n337), .A2(new_n338), .A3(new_n332), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n329), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  XNOR2_X1  g139(.A(G113gat), .B(G120gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(KEYINPUT70), .ZN(new_n342));
  INV_X1    g141(.A(G134gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(G127gat), .ZN(new_n344));
  INV_X1    g143(.A(G127gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G134gat), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n344), .A2(new_n346), .A3(new_n331), .ZN(new_n347));
  NAND4_X1  g146(.A1(new_n342), .A2(new_n347), .A3(KEYINPUT71), .A4(new_n334), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n331), .B1(new_n337), .B2(new_n338), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT69), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n351), .B1(new_n350), .B2(new_n330), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n340), .A2(new_n348), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(G141gat), .ZN(new_n354));
  INV_X1    g153(.A(G148gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(G141gat), .A2(G148gat), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n356), .A2(KEYINPUT81), .A3(new_n357), .ZN(new_n361));
  NAND2_X1  g160(.A1(G155gat), .A2(G162gat), .ZN(new_n362));
  OR3_X1    g161(.A1(KEYINPUT2), .A2(G155gat), .A3(G162gat), .ZN(new_n363));
  AOI22_X1  g162(.A1(new_n360), .A2(new_n361), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT80), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g165(.A1(KEYINPUT80), .A2(G155gat), .A3(G162gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n366), .B(new_n367), .C1(KEYINPUT79), .C2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n358), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n362), .A2(KEYINPUT2), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n366), .A2(new_n367), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n368), .A2(KEYINPUT79), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n370), .A2(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n364), .B1(new_n369), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n353), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n370), .A2(new_n371), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n372), .A2(new_n373), .ZN(new_n380));
  AND3_X1   g179(.A1(new_n379), .A2(new_n380), .A3(new_n369), .ZN(new_n381));
  OAI21_X1  g180(.A(KEYINPUT3), .B1(new_n381), .B2(new_n364), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n340), .A2(new_n348), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n352), .A2(new_n349), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n364), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n374), .A2(new_n369), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT3), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n382), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n353), .A2(new_n375), .A3(KEYINPUT4), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n378), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(G225gat), .A2(G233gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  AND2_X1   g193(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT39), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n328), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n387), .A2(new_n386), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n385), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT82), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n400), .A3(new_n376), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n385), .A2(KEYINPUT82), .A3(new_n398), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n394), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OR2_X1    g202(.A1(new_n395), .A2(new_n396), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n397), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT40), .ZN(new_n406));
  OR2_X1    g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n401), .A2(new_n394), .A3(new_n402), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(KEYINPUT5), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n378), .A2(new_n390), .A3(new_n393), .A4(new_n391), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT5), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(new_n328), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n405), .A2(new_n406), .ZN(new_n416));
  AND3_X1   g215(.A1(new_n407), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n316), .A2(new_n323), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(G228gat), .A2(G233gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n389), .A2(new_n263), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n419), .B1(new_n420), .B2(new_n281), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n388), .B1(new_n281), .B2(KEYINPUT29), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n398), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n388), .B1(new_n281), .B2(new_n264), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n398), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n420), .A2(new_n281), .ZN(new_n428));
  AOI22_X1  g227(.A1(new_n427), .A2(new_n428), .B1(G228gat), .B2(G233gat), .ZN(new_n429));
  OAI21_X1  g228(.A(G22gat), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT87), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G78gat), .B(G106gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(G50gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n434), .B(KEYINPUT86), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n435), .B(KEYINPUT31), .Z(new_n436));
  INV_X1    g235(.A(new_n429), .ZN(new_n437));
  INV_X1    g236(.A(G22gat), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n438), .A3(new_n424), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n432), .A2(new_n436), .B1(new_n439), .B2(new_n430), .ZN(new_n440));
  AND4_X1   g239(.A1(KEYINPUT87), .A2(new_n439), .A3(new_n430), .A4(new_n436), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(KEYINPUT89), .B(KEYINPUT37), .Z(new_n444));
  NAND2_X1  g243(.A1(new_n282), .A2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n446), .B1(new_n303), .B2(new_n304), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT37), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n447), .B(new_n321), .C1(new_n312), .C2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT38), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n411), .A2(KEYINPUT6), .A3(new_n328), .A4(new_n414), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT85), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n413), .B1(new_n409), .B2(new_n410), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT85), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT6), .A4(new_n328), .ZN(new_n455));
  AND2_X1   g254(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n411), .A2(new_n414), .ZN(new_n457));
  INV_X1    g256(.A(new_n328), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT6), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n460), .A3(new_n415), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n317), .A2(new_n456), .A3(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT38), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n448), .B1(new_n274), .B2(new_n300), .ZN(new_n465));
  INV_X1    g264(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n299), .A2(new_n281), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n467), .B1(new_n294), .B2(new_n297), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n464), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n447), .A2(new_n470), .A3(new_n321), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT90), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n310), .A2(new_n311), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n285), .B1(new_n474), .B2(new_n446), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n475), .A2(KEYINPUT90), .A3(new_n470), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n450), .A2(new_n463), .A3(new_n473), .A4(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n418), .A2(new_n443), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT84), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n415), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n453), .A2(KEYINPUT84), .A3(new_n328), .ZN(new_n481));
  NAND4_X1  g280(.A1(new_n480), .A2(new_n459), .A3(new_n460), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n456), .A2(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n319), .A2(new_n483), .A3(new_n322), .A4(new_n305), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n442), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n290), .A2(new_n353), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n260), .A2(new_n385), .ZN(new_n487));
  INV_X1    g286(.A(G227gat), .ZN(new_n488));
  INV_X1    g287(.A(G233gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n486), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT32), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT72), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n491), .A2(KEYINPUT72), .A3(KEYINPUT32), .ZN(new_n495));
  XNOR2_X1  g294(.A(G15gat), .B(G43gat), .ZN(new_n496));
  XNOR2_X1  g295(.A(G71gat), .B(G99gat), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n496), .B(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT33), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(new_n491), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n494), .A2(new_n495), .A3(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n491), .B(KEYINPUT32), .C1(new_n499), .C2(new_n498), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT34), .ZN(new_n504));
  INV_X1    g303(.A(new_n490), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n504), .B1(new_n503), .B2(new_n505), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n501), .A2(new_n502), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n509), .B1(new_n501), .B2(new_n502), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT36), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT36), .ZN(new_n515));
  OAI21_X1  g314(.A(new_n515), .B1(new_n511), .B2(new_n512), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n485), .A2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n316), .A2(new_n323), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT91), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n521), .B1(new_n511), .B2(new_n512), .ZN(new_n522));
  INV_X1    g321(.A(new_n512), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(KEYINPUT91), .A3(new_n510), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  AOI211_X1 g324(.A(KEYINPUT35), .B(new_n442), .C1(new_n456), .C2(new_n461), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n520), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n313), .A2(new_n315), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n442), .A2(new_n511), .A3(new_n512), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(new_n483), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT35), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n478), .A2(new_n519), .B1(new_n527), .B2(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(G113gat), .B(G141gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n533), .B(G197gat), .ZN(new_n534));
  XOR2_X1   g333(.A(KEYINPUT11), .B(G169gat), .Z(new_n535));
  XNOR2_X1  g334(.A(new_n534), .B(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n536), .B(KEYINPUT12), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(G15gat), .B(G22gat), .ZN(new_n539));
  INV_X1    g338(.A(G1gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n540), .A2(KEYINPUT93), .A3(KEYINPUT16), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT93), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT16), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(G1gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(new_n541), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(G1gat), .B2(new_n539), .ZN(new_n546));
  OAI21_X1  g345(.A(KEYINPUT94), .B1(new_n539), .B2(G1gat), .ZN(new_n547));
  INV_X1    g346(.A(G8gat), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n546), .B(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(G29gat), .A2(G36gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT14), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G29gat), .ZN(new_n554));
  INV_X1    g353(.A(G36gat), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(G43gat), .B(G50gat), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n557), .A2(KEYINPUT15), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT92), .B1(new_n554), .B2(new_n555), .ZN(new_n560));
  OR3_X1    g359(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT92), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n553), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  XNOR2_X1  g361(.A(new_n557), .B(KEYINPUT15), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n559), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AND2_X1   g363(.A1(new_n550), .A2(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(KEYINPUT17), .ZN(new_n566));
  INV_X1    g365(.A(new_n550), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G229gat), .A2(G233gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT95), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(KEYINPUT18), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n568), .A2(new_n569), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n550), .B(new_n564), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n569), .B(KEYINPUT13), .Z(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n572), .B1(new_n568), .B2(new_n569), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n538), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n578), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n580), .A2(new_n537), .A3(new_n576), .A4(new_n573), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n532), .A2(new_n583), .ZN(new_n584));
  AND2_X1   g383(.A1(G232gat), .A2(G233gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n585), .A2(KEYINPUT41), .ZN(new_n586));
  XNOR2_X1  g385(.A(G134gat), .B(G162gat), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT102), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n590), .B(KEYINPUT103), .Z(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G85gat), .A2(G92gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT7), .ZN(new_n594));
  NAND2_X1  g393(.A1(G99gat), .A2(G106gat), .ZN(new_n595));
  INV_X1    g394(.A(G85gat), .ZN(new_n596));
  INV_X1    g395(.A(G92gat), .ZN(new_n597));
  AOI22_X1  g396(.A1(KEYINPUT8), .A2(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n594), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G99gat), .B(G106gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  NAND2_X1  g400(.A1(new_n566), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n599), .B(new_n600), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n564), .A2(new_n603), .B1(KEYINPUT41), .B2(new_n585), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT101), .ZN(new_n606));
  XNOR2_X1  g405(.A(G190gat), .B(G218gat), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT101), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n602), .A2(new_n608), .A3(new_n604), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n606), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  OR2_X1    g409(.A1(new_n588), .A2(new_n589), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI21_X1  g411(.A(new_n607), .B1(new_n606), .B2(new_n609), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n592), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n613), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n615), .A2(new_n611), .A3(new_n610), .A4(new_n591), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT98), .ZN(new_n618));
  XOR2_X1   g417(.A(G57gat), .B(G64gat), .Z(new_n619));
  NAND2_X1  g418(.A1(G71gat), .A2(G78gat), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT9), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n622), .A2(KEYINPUT97), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT97), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n620), .A2(new_n624), .A3(new_n621), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n619), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g425(.A(G71gat), .B(G78gat), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(KEYINPUT96), .A3(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n627), .B1(new_n626), .B2(KEYINPUT96), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n618), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n626), .A2(KEYINPUT96), .ZN(new_n632));
  INV_X1    g431(.A(new_n627), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n634), .A2(KEYINPUT98), .A3(new_n628), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n637), .A2(KEYINPUT21), .ZN(new_n638));
  INV_X1    g437(.A(G231gat), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n639), .A2(new_n489), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n638), .A2(new_n641), .ZN(new_n644));
  OAI21_X1  g443(.A(G127gat), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n644), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n646), .A2(new_n345), .A3(new_n642), .ZN(new_n647));
  XNOR2_X1  g446(.A(G183gat), .B(G211gat), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n645), .A2(new_n647), .A3(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n649), .B1(new_n645), .B2(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n637), .A2(KEYINPUT21), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT99), .B(KEYINPUT100), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n653), .A2(new_n567), .A3(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n654), .B1(new_n653), .B2(new_n567), .ZN(new_n656));
  XNOR2_X1  g455(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n657));
  INV_X1    g456(.A(G155gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  OR3_X1    g458(.A1(new_n655), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n659), .B1(new_n655), .B2(new_n656), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OR3_X1    g461(.A1(new_n651), .A2(new_n652), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n662), .B1(new_n651), .B2(new_n652), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n617), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(G230gat), .A2(G233gat), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n631), .A2(new_n601), .A3(new_n635), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n603), .A2(new_n634), .A3(new_n628), .ZN(new_n669));
  AOI21_X1  g468(.A(KEYINPUT10), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND4_X1   g469(.A1(KEYINPUT10), .A2(new_n631), .A3(new_n635), .A4(new_n603), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n667), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n668), .A2(G230gat), .A3(G233gat), .A4(new_n669), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(G120gat), .B(G148gat), .ZN(new_n675));
  XNOR2_X1  g474(.A(G176gat), .B(G204gat), .ZN(new_n676));
  XOR2_X1   g475(.A(new_n675), .B(new_n676), .Z(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n672), .A2(new_n673), .A3(new_n677), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n584), .A2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n483), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(new_n540), .ZN(G1324gat));
  NOR3_X1   g484(.A1(new_n520), .A2(new_n666), .A3(new_n681), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT16), .B(G8gat), .Z(new_n687));
  AND3_X1   g486(.A1(new_n584), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n548), .B1(new_n584), .B2(new_n686), .ZN(new_n689));
  OAI21_X1  g488(.A(KEYINPUT42), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n690), .B1(KEYINPUT42), .B2(new_n688), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT104), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693));
  OAI211_X1 g492(.A(new_n690), .B(new_n693), .C1(KEYINPUT42), .C2(new_n688), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(G1325gat));
  OAI21_X1  g494(.A(G15gat), .B1(new_n683), .B2(new_n517), .ZN(new_n696));
  INV_X1    g495(.A(G15gat), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n584), .A2(new_n697), .A3(new_n525), .A4(new_n682), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT105), .ZN(G1326gat));
  NOR2_X1   g499(.A1(new_n683), .A2(new_n443), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT43), .B(G22gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1327gat));
  AOI21_X1  g502(.A(KEYINPUT90), .B1(new_n475), .B2(new_n470), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n445), .B1(new_n310), .B2(new_n311), .ZN(new_n705));
  NOR4_X1   g504(.A1(new_n705), .A2(new_n469), .A3(new_n472), .A4(new_n285), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n462), .B1(new_n449), .B2(KEYINPUT38), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n442), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n518), .B1(new_n709), .B2(new_n418), .ZN(new_n710));
  INV_X1    g509(.A(new_n525), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n711), .B1(new_n316), .B2(new_n323), .ZN(new_n712));
  AOI22_X1  g511(.A1(new_n712), .A2(new_n526), .B1(new_n530), .B2(KEYINPUT35), .ZN(new_n713));
  OAI21_X1  g512(.A(KEYINPUT107), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n478), .A2(new_n519), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n527), .A2(new_n531), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n617), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n719), .A2(KEYINPUT44), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n714), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(KEYINPUT44), .B1(new_n532), .B2(new_n719), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AND3_X1   g522(.A1(new_n664), .A2(KEYINPUT106), .A3(new_n663), .ZN(new_n724));
  AOI21_X1  g523(.A(KEYINPUT106), .B1(new_n663), .B2(new_n664), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n727), .A2(new_n583), .A3(new_n681), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n723), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(G29gat), .B1(new_n729), .B2(new_n483), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT45), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n715), .A2(new_n717), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n663), .A2(new_n664), .ZN(new_n733));
  NOR3_X1   g532(.A1(new_n733), .A2(new_n719), .A3(new_n681), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n732), .A2(new_n582), .A3(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n483), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n554), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n731), .B1(new_n735), .B2(new_n737), .ZN(new_n738));
  OR3_X1    g537(.A1(new_n735), .A2(new_n731), .A3(new_n737), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n730), .A2(new_n738), .A3(new_n739), .ZN(G1328gat));
  OAI21_X1  g539(.A(G36gat), .B1(new_n729), .B2(new_n520), .ZN(new_n741));
  INV_X1    g540(.A(new_n520), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(new_n555), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT46), .B1(new_n735), .B2(new_n743), .ZN(new_n744));
  OR3_X1    g543(.A1(new_n735), .A2(KEYINPUT46), .A3(new_n743), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n741), .A2(new_n744), .A3(new_n745), .ZN(G1329gat));
  XNOR2_X1  g545(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n747));
  INV_X1    g546(.A(new_n517), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n723), .A2(new_n748), .A3(new_n728), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(G43gat), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n735), .A2(G43gat), .A3(new_n711), .ZN(new_n751));
  INV_X1    g550(.A(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n747), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n747), .ZN(new_n754));
  AOI211_X1 g553(.A(new_n751), .B(new_n754), .C1(new_n749), .C2(G43gat), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n753), .A2(new_n755), .ZN(G1330gat));
  NAND3_X1  g555(.A1(new_n723), .A2(new_n442), .A3(new_n728), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n757), .A2(G50gat), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT110), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n443), .A2(G50gat), .ZN(new_n760));
  INV_X1    g559(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n759), .B1(new_n735), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n584), .A2(KEYINPUT110), .A3(new_n734), .A4(new_n760), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n762), .A2(KEYINPUT48), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT109), .B1(new_n735), .B2(new_n761), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n584), .A2(new_n766), .A3(new_n734), .A4(new_n760), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n768), .B1(new_n757), .B2(G50gat), .ZN(new_n769));
  OAI22_X1  g568(.A1(new_n758), .A2(new_n764), .B1(new_n769), .B2(KEYINPUT48), .ZN(G1331gat));
  AND2_X1   g569(.A1(new_n714), .A2(new_n718), .ZN(new_n771));
  INV_X1    g570(.A(new_n681), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n666), .A2(new_n582), .A3(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(new_n736), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n742), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n778), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n779));
  XOR2_X1   g578(.A(KEYINPUT49), .B(G64gat), .Z(new_n780));
  OAI21_X1  g579(.A(new_n779), .B1(new_n778), .B2(new_n780), .ZN(G1333gat));
  NAND4_X1  g580(.A1(new_n714), .A2(new_n718), .A3(new_n748), .A4(new_n773), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(G71gat), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n711), .A2(G71gat), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n783), .B1(new_n774), .B2(new_n784), .ZN(new_n785));
  XOR2_X1   g584(.A(new_n785), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g585(.A1(new_n775), .A2(new_n442), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g587(.A1(new_n483), .A2(G85gat), .A3(new_n772), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n733), .A2(new_n582), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n732), .A2(new_n617), .A3(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n732), .A2(KEYINPUT51), .A3(new_n617), .A4(new_n790), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n793), .A2(KEYINPUT112), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(KEYINPUT112), .B1(new_n793), .B2(new_n794), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n789), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n790), .A2(new_n681), .ZN(new_n798));
  INV_X1    g597(.A(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n723), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT111), .B1(new_n800), .B2(new_n483), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G85gat), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n800), .A2(KEYINPUT111), .A3(new_n483), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n797), .B1(new_n802), .B2(new_n803), .ZN(G1336gat));
  AND3_X1   g603(.A1(new_n791), .A2(KEYINPUT114), .A3(KEYINPUT51), .ZN(new_n805));
  AOI21_X1  g604(.A(KEYINPUT51), .B1(new_n791), .B2(KEYINPUT114), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n742), .A2(new_n597), .A3(new_n681), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n807), .B(KEYINPUT113), .ZN(new_n808));
  NOR3_X1   g607(.A1(new_n805), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  AOI21_X1  g608(.A(new_n798), .B1(new_n721), .B2(new_n722), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n597), .B1(new_n810), .B2(new_n742), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n793), .A2(new_n794), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(new_n808), .ZN(new_n815));
  OAI22_X1  g614(.A1(new_n812), .A2(new_n813), .B1(new_n811), .B2(new_n815), .ZN(G1337gat));
  NOR3_X1   g615(.A1(new_n711), .A2(G99gat), .A3(new_n772), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n817), .B(KEYINPUT115), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n795), .B2(new_n796), .ZN(new_n819));
  OAI21_X1  g618(.A(G99gat), .B1(new_n800), .B2(new_n517), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(G1338gat));
  NOR3_X1   g620(.A1(new_n443), .A2(G106gat), .A3(new_n772), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n805), .A2(new_n806), .A3(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(G106gat), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n810), .B2(new_n442), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n828), .B1(new_n814), .B2(new_n823), .ZN(new_n829));
  OAI22_X1  g628(.A1(new_n827), .A2(new_n828), .B1(new_n826), .B2(new_n829), .ZN(G1339gat));
  NAND3_X1  g629(.A1(new_n665), .A2(new_n583), .A3(new_n772), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT116), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n665), .A2(new_n833), .A3(new_n583), .A4(new_n772), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836));
  OAI211_X1 g635(.A(new_n836), .B(new_n667), .C1(new_n670), .C2(new_n671), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n678), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n672), .A2(KEYINPUT54), .ZN(new_n839));
  OR3_X1    g638(.A1(new_n670), .A2(new_n667), .A3(new_n671), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(KEYINPUT55), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n680), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT117), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n839), .A2(new_n840), .ZN(new_n845));
  INV_X1    g644(.A(new_n838), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT55), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n843), .A2(KEYINPUT117), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n844), .A2(new_n582), .A3(new_n849), .A4(new_n850), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n568), .A2(new_n569), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n574), .A2(new_n575), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n536), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n581), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n681), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n617), .B1(new_n851), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n855), .A2(new_n614), .A3(new_n616), .ZN(new_n858));
  AND4_X1   g657(.A1(new_n844), .A2(new_n858), .A3(new_n849), .A4(new_n850), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n726), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n835), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n483), .A2(new_n442), .ZN(new_n862));
  AND4_X1   g661(.A1(new_n520), .A2(new_n861), .A3(new_n513), .A4(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(G113gat), .B1(new_n863), .B2(new_n582), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n861), .A2(new_n712), .A3(new_n862), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n583), .A2(new_n336), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(G1340gat));
  AOI21_X1  g666(.A(G120gat), .B1(new_n863), .B2(new_n681), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n772), .A2(new_n333), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n868), .B1(new_n865), .B2(new_n869), .ZN(G1341gat));
  NAND3_X1  g669(.A1(new_n865), .A2(G127gat), .A3(new_n727), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(KEYINPUT118), .ZN(new_n873));
  AOI21_X1  g672(.A(G127gat), .B1(new_n863), .B2(new_n733), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G1342gat));
  NAND3_X1  g674(.A1(new_n863), .A2(new_n343), .A3(new_n617), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(KEYINPUT56), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n343), .B1(new_n865), .B2(new_n617), .ZN(new_n879));
  OR3_X1    g678(.A1(new_n877), .A2(new_n878), .A3(new_n879), .ZN(G1343gat));
  INV_X1    g679(.A(KEYINPUT121), .ZN(new_n881));
  INV_X1    g680(.A(new_n733), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n847), .A2(KEYINPUT119), .A3(new_n848), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n884), .B1(new_n841), .B2(KEYINPUT55), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n582), .A2(new_n842), .A3(new_n680), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n856), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n617), .B1(new_n888), .B2(new_n889), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n881), .B(new_n882), .C1(new_n892), .C2(new_n859), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n859), .B1(new_n890), .B2(new_n891), .ZN(new_n894));
  OAI21_X1  g693(.A(KEYINPUT121), .B1(new_n894), .B2(new_n733), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n893), .A2(new_n895), .A3(new_n835), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT57), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n443), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n861), .A2(new_n442), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n897), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n742), .A2(new_n483), .A3(new_n748), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n902), .A2(new_n582), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(G141gat), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n906));
  INV_X1    g705(.A(new_n903), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n900), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n908), .A2(new_n354), .A3(new_n582), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n905), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n907), .B1(new_n899), .B2(new_n901), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n354), .B1(new_n911), .B2(new_n582), .ZN(new_n912));
  INV_X1    g711(.A(new_n909), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT58), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n910), .A2(new_n914), .ZN(G1344gat));
  NAND3_X1  g714(.A1(new_n908), .A2(new_n355), .A3(new_n681), .ZN(new_n916));
  AOI211_X1 g715(.A(KEYINPUT59), .B(new_n355), .C1(new_n911), .C2(new_n681), .ZN(new_n917));
  XNOR2_X1  g716(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n900), .A2(new_n897), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n831), .B1(new_n894), .B2(new_n733), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT57), .B1(new_n920), .B2(new_n442), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n681), .B(new_n903), .C1(new_n919), .C2(new_n921), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n918), .B1(new_n922), .B2(G148gat), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n916), .B1(new_n917), .B2(new_n923), .ZN(G1345gat));
  INV_X1    g723(.A(new_n911), .ZN(new_n925));
  OAI21_X1  g724(.A(G155gat), .B1(new_n925), .B2(new_n726), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n908), .A2(new_n658), .A3(new_n733), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(G1346gat));
  OAI21_X1  g727(.A(G162gat), .B1(new_n925), .B2(new_n719), .ZN(new_n929));
  INV_X1    g728(.A(G162gat), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n908), .A2(new_n930), .A3(new_n617), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n929), .A2(new_n931), .ZN(G1347gat));
  NOR2_X1   g731(.A1(new_n520), .A2(new_n736), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n711), .A2(new_n442), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n861), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n861), .A2(new_n933), .A3(KEYINPUT123), .A4(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(G169gat), .B1(new_n939), .B2(new_n583), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n861), .A2(new_n529), .A3(new_n933), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n941), .A2(new_n229), .A3(new_n230), .A4(new_n582), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(G1348gat));
  OAI21_X1  g742(.A(G176gat), .B1(new_n939), .B2(new_n772), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n941), .A2(new_n216), .A3(new_n681), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1349gat));
  OAI21_X1  g745(.A(G183gat), .B1(new_n939), .B2(new_n726), .ZN(new_n947));
  AND2_X1   g746(.A1(new_n733), .A2(new_n211), .ZN(new_n948));
  AOI21_X1  g747(.A(KEYINPUT124), .B1(new_n941), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(KEYINPUT60), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT60), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n947), .A2(new_n952), .A3(new_n949), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n951), .A2(new_n953), .ZN(G1350gat));
  NAND3_X1  g753(.A1(new_n941), .A2(new_n207), .A3(new_n617), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n937), .A2(new_n617), .A3(new_n938), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  AND4_X1   g756(.A1(KEYINPUT125), .A2(new_n956), .A3(new_n957), .A4(G190gat), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n207), .B1(new_n959), .B2(KEYINPUT61), .ZN(new_n960));
  AOI22_X1  g759(.A1(new_n956), .A2(new_n960), .B1(KEYINPUT125), .B2(new_n957), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n955), .B1(new_n958), .B2(new_n961), .ZN(G1351gat));
  NAND2_X1  g761(.A1(new_n933), .A2(new_n517), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n900), .A2(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(G197gat), .B1(new_n964), .B2(new_n582), .ZN(new_n965));
  OR2_X1    g764(.A1(new_n919), .A2(new_n921), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n963), .B(KEYINPUT126), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n582), .A2(G197gat), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(G1352gat));
  NAND3_X1  g769(.A1(new_n966), .A2(new_n681), .A3(new_n967), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n971), .A2(G204gat), .ZN(new_n972));
  NOR4_X1   g771(.A1(new_n900), .A2(G204gat), .A3(new_n772), .A4(new_n963), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT62), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(G1353gat));
  INV_X1    g774(.A(G211gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n964), .A2(new_n976), .A3(new_n733), .ZN(new_n977));
  OAI211_X1 g776(.A(new_n967), .B(new_n733), .C1(new_n919), .C2(new_n921), .ZN(new_n978));
  AND3_X1   g777(.A1(new_n978), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n979));
  AOI21_X1  g778(.A(KEYINPUT63), .B1(new_n978), .B2(G211gat), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n977), .B1(new_n979), .B2(new_n980), .ZN(G1354gat));
  AOI21_X1  g780(.A(G218gat), .B1(new_n964), .B2(new_n617), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n617), .A2(G218gat), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT127), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n982), .B1(new_n968), .B2(new_n984), .ZN(G1355gat));
endmodule


