//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:06 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1262, new_n1263,
    new_n1264;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0005(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n206));
  INV_X1    g0006(.A(G116), .ZN(new_n207));
  INV_X1    g0007(.A(G270), .ZN(new_n208));
  OAI21_X1  g0008(.A(new_n206), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G68), .A2(G238), .ZN(new_n211));
  INV_X1    g0011(.A(G50), .ZN(new_n212));
  INV_X1    g0012(.A(G226), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n210), .B(new_n211), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n214), .C1(G97), .C2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G1), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT1), .Z(new_n220));
  NAND2_X1  g0020(.A1(new_n203), .A2(G50), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT65), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n223), .A2(new_n217), .A3(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(KEYINPUT64), .ZN(new_n226));
  INV_X1    g0026(.A(new_n218), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n226), .B1(new_n227), .B2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G13), .ZN(new_n229));
  NAND3_X1  g0029(.A1(new_n218), .A2(KEYINPUT64), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n231), .B(G250), .C1(G257), .C2(G264), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(KEYINPUT0), .Z(new_n233));
  NOR3_X1   g0033(.A1(new_n220), .A2(new_n225), .A3(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G226), .B(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(G238), .B(G244), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n224), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n217), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n217), .A2(new_n256), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n253), .A2(new_n254), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n258), .B(KEYINPUT70), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n203), .A2(G50), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n217), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n252), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n216), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(new_n252), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n216), .A2(G20), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n265), .A2(G50), .A3(new_n266), .ZN(new_n267));
  AND2_X1   g0067(.A1(new_n262), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n268), .B1(G50), .B2(new_n263), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n268), .B(KEYINPUT9), .C1(G50), .C2(new_n263), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G274), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT67), .B(G45), .ZN(new_n275));
  INV_X1    g0075(.A(G41), .ZN(new_n276));
  AOI21_X1  g0076(.A(G1), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT68), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT67), .A2(G45), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT67), .A2(G45), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n276), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(new_n216), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n280), .B1(new_n284), .B2(KEYINPUT68), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  AOI21_X1  g0087(.A(G1), .B1(new_n276), .B2(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n280), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(G226), .ZN(new_n290));
  XNOR2_X1  g0090(.A(KEYINPUT3), .B(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G223), .A2(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G222), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n291), .A2(new_n292), .A3(new_n294), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n295), .B(new_n280), .C1(G77), .C2(new_n291), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n286), .A2(new_n290), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g0097(.A(new_n297), .B(KEYINPUT69), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(G200), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(G190), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT72), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n273), .B(new_n302), .C1(new_n303), .C2(KEYINPUT10), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n271), .A2(new_n300), .A3(new_n301), .A4(new_n272), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n300), .A2(new_n303), .A3(new_n301), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G179), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n298), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n310), .B(new_n269), .C1(G169), .C2(new_n298), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n304), .A2(new_n308), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n289), .A2(G244), .ZN(new_n313));
  NAND2_X1  g0113(.A1(G238), .A2(G1698), .ZN(new_n314));
  INV_X1    g0114(.A(G232), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n291), .B(new_n314), .C1(new_n315), .C2(G1698), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n316), .B(new_n280), .C1(G107), .C2(new_n291), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n286), .A2(new_n313), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(G169), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n319), .B1(new_n309), .B2(new_n318), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n263), .B(KEYINPUT71), .ZN(new_n321));
  INV_X1    g0121(.A(G77), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n321), .ZN(new_n324));
  INV_X1    g0124(.A(new_n252), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n324), .A2(new_n325), .A3(new_n266), .ZN(new_n326));
  XOR2_X1   g0126(.A(KEYINPUT15), .B(G87), .Z(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n253), .A2(new_n257), .B1(new_n328), .B2(new_n254), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(G20), .B2(G77), .ZN(new_n330));
  OAI221_X1 g0130(.A(new_n323), .B1(new_n322), .B2(new_n326), .C1(new_n330), .C2(new_n325), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n320), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n318), .A2(G200), .ZN(new_n333));
  INV_X1    g0133(.A(G190), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n334), .B2(new_n318), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n332), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n326), .A2(new_n202), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n202), .A2(G20), .ZN(new_n338));
  OAI221_X1 g0138(.A(new_n338), .B1(new_n254), .B2(new_n322), .C1(new_n212), .C2(new_n257), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n252), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT11), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT12), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n321), .B2(new_n202), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT74), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n344), .B(new_n345), .ZN(new_n346));
  NOR4_X1   g0146(.A1(new_n338), .A2(KEYINPUT12), .A3(G1), .A4(new_n229), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AOI211_X1 g0148(.A(new_n337), .B(new_n342), .C1(new_n346), .C2(new_n348), .ZN(new_n349));
  AOI22_X1  g0149(.A1(new_n279), .A2(new_n285), .B1(G238), .B2(new_n289), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT73), .ZN(new_n351));
  INV_X1    g0151(.A(G97), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n256), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g0153(.A1(G226), .A2(G1698), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n354), .B1(new_n315), .B2(G1698), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n353), .B1(new_n355), .B2(new_n291), .ZN(new_n356));
  INV_X1    g0156(.A(new_n224), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(new_n256), .B2(new_n276), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n351), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n315), .A2(G1698), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(G226), .B2(G1698), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT3), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(G33), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g0166(.A(KEYINPUT73), .B(new_n280), .C1(new_n366), .C2(new_n353), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n359), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  AND3_X1   g0169(.A1(new_n350), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n369), .B1(new_n350), .B2(new_n368), .ZN(new_n371));
  OAI21_X1  g0171(.A(G200), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n371), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n350), .A2(new_n369), .A3(new_n368), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(G190), .A3(new_n374), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n349), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n370), .A2(new_n371), .ZN(new_n377));
  INV_X1    g0177(.A(G169), .ZN(new_n378));
  OAI21_X1  g0178(.A(KEYINPUT14), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(G179), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT14), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(G169), .C1(new_n370), .C2(new_n371), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(new_n349), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n376), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT77), .ZN(new_n387));
  XNOR2_X1  g0187(.A(G58), .B(G68), .ZN(new_n388));
  INV_X1    g0188(.A(new_n257), .ZN(new_n389));
  AOI22_X1  g0189(.A1(G20), .A2(new_n388), .B1(new_n389), .B2(G159), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n363), .A2(G33), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n256), .A2(KEYINPUT3), .ZN(new_n392));
  OAI211_X1 g0192(.A(KEYINPUT7), .B(new_n217), .C1(new_n391), .C2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n362), .A2(new_n364), .A3(KEYINPUT75), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT75), .B1(new_n362), .B2(new_n364), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n217), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  OAI211_X1 g0199(.A(KEYINPUT16), .B(new_n390), .C1(new_n399), .C2(new_n202), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n252), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT76), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n393), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n398), .B1(new_n291), .B2(G20), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n365), .A2(KEYINPUT76), .A3(KEYINPUT7), .A4(new_n217), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(G68), .ZN(new_n407));
  AOI21_X1  g0207(.A(KEYINPUT16), .B1(new_n407), .B2(new_n390), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n387), .B1(new_n401), .B2(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n253), .B1(new_n216), .B2(G20), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n410), .A2(new_n265), .B1(new_n264), .B2(new_n253), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n407), .A2(new_n390), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT16), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n414), .A2(KEYINPUT77), .A3(new_n252), .A4(new_n400), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n409), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n362), .A2(new_n364), .A3(G223), .A4(new_n293), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT78), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n291), .A2(KEYINPUT78), .A3(G223), .A4(new_n293), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G87), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n291), .A2(G226), .A3(G1698), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n419), .A2(new_n420), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n280), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n289), .A2(G232), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n424), .A2(new_n286), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(G169), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n424), .A2(new_n286), .A3(G179), .A4(new_n425), .ZN(new_n428));
  AOI21_X1  g0228(.A(KEYINPUT79), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n427), .A2(KEYINPUT79), .A3(new_n428), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT18), .B1(new_n416), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(G200), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n426), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g0235(.A(new_n435), .B1(G190), .B2(new_n426), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n416), .A2(KEYINPUT17), .A3(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n409), .A2(new_n415), .A3(new_n411), .A4(new_n436), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT17), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n427), .A2(KEYINPUT79), .A3(new_n428), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(new_n429), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n409), .A2(new_n415), .A3(new_n411), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT18), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  NAND4_X1  g0245(.A1(new_n433), .A2(new_n437), .A3(new_n440), .A4(new_n445), .ZN(new_n446));
  NOR4_X1   g0246(.A1(new_n312), .A2(new_n336), .A3(new_n386), .A4(new_n446), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n362), .A2(new_n364), .A3(new_n217), .A4(G87), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT22), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT22), .ZN(new_n450));
  NAND4_X1  g0250(.A1(new_n291), .A2(new_n450), .A3(new_n217), .A4(G87), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n256), .A2(new_n207), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n217), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n217), .A2(G107), .ZN(new_n455));
  XNOR2_X1  g0255(.A(new_n455), .B(KEYINPUT23), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n452), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT24), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n449), .A2(new_n451), .B1(new_n217), .B2(new_n453), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT24), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n459), .A2(new_n460), .A3(new_n456), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n325), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n216), .A2(G33), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n265), .A2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(G107), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT87), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n467), .A2(KEYINPUT25), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n263), .A2(new_n468), .A3(G107), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n467), .A2(KEYINPUT25), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n469), .B(new_n470), .ZN(new_n471));
  NOR3_X1   g0271(.A1(new_n462), .A2(new_n466), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(G257), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(G1698), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n291), .B(new_n474), .C1(G250), .C2(G1698), .ZN(new_n475));
  NAND2_X1  g0275(.A1(G33), .A2(G294), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(new_n280), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n287), .A2(G1), .ZN(new_n479));
  AND2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  NOR2_X1   g0280(.A1(KEYINPUT5), .A2(G41), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  OR2_X1    g0282(.A1(new_n482), .A2(new_n274), .ZN(new_n483));
  AND2_X1   g0283(.A1(new_n482), .A2(new_n358), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(G264), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n478), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(new_n334), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n486), .A2(G200), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n472), .A2(new_n488), .A3(KEYINPUT89), .A4(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT89), .ZN(new_n491));
  AND4_X1   g0291(.A1(new_n460), .A2(new_n452), .A3(new_n454), .A4(new_n456), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n460), .B1(new_n459), .B2(new_n456), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n252), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n466), .ZN(new_n495));
  INV_X1    g0295(.A(new_n471), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n494), .A2(new_n489), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n491), .B1(new_n497), .B2(new_n487), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n490), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n263), .A2(G97), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n406), .A2(G107), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n465), .A2(KEYINPUT6), .A3(G97), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n352), .A2(new_n465), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G97), .A2(G107), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n502), .B1(new_n505), .B2(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G20), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n389), .A2(G77), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n501), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n500), .B1(new_n509), .B2(new_n252), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n464), .A2(new_n352), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n362), .A2(new_n364), .A3(G244), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT4), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G283), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n514), .A2(G1698), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n517), .A2(new_n362), .A3(new_n364), .A4(G244), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n362), .A2(new_n364), .A3(G250), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n293), .B1(new_n520), .B2(KEYINPUT4), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n280), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n484), .A2(G257), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n483), .A3(new_n523), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n524), .A2(KEYINPUT80), .A3(G200), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT80), .B1(new_n524), .B2(G200), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n510), .B(new_n512), .C1(new_n525), .C2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n522), .A2(G190), .A3(new_n483), .A4(new_n523), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT81), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n528), .B(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(KEYINPUT82), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n510), .A2(new_n512), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n524), .A2(new_n378), .ZN(new_n533));
  INV_X1    g0333(.A(new_n524), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n309), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n526), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n524), .A2(KEYINPUT80), .A3(G200), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n528), .B(KEYINPUT81), .ZN(new_n540));
  AOI211_X1 g0340(.A(new_n500), .B(new_n511), .C1(new_n509), .C2(new_n252), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT82), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n539), .A2(new_n540), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  AND4_X1   g0343(.A1(new_n499), .A2(new_n531), .A3(new_n536), .A4(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n516), .B(new_n217), .C1(G33), .C2(new_n352), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n545), .B(new_n252), .C1(new_n217), .C2(G116), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT20), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n546), .B1(KEYINPUT85), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(KEYINPUT85), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  OR2_X1    g0350(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n321), .A2(new_n207), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n550), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n324), .A2(G116), .A3(new_n325), .A4(new_n463), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n551), .A2(new_n552), .A3(new_n553), .A4(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n484), .A2(G270), .ZN(new_n557));
  INV_X1    g0357(.A(G303), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n358), .B1(new_n558), .B2(new_n365), .ZN(new_n559));
  NAND2_X1  g0359(.A1(G264), .A2(G1698), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n291), .B(new_n560), .C1(new_n473), .C2(G1698), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n559), .A2(KEYINPUT84), .A3(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g0363(.A(KEYINPUT84), .B1(new_n559), .B2(new_n561), .ZN(new_n564));
  OAI211_X1 g0364(.A(new_n483), .B(new_n557), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(G200), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n556), .B(new_n566), .C1(new_n334), .C2(new_n565), .ZN(new_n567));
  INV_X1    g0367(.A(new_n479), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n358), .A2(G250), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n479), .A2(G274), .ZN(new_n570));
  MUX2_X1   g0370(.A(G238), .B(G244), .S(G1698), .Z(new_n571));
  AOI21_X1  g0371(.A(new_n453), .B1(new_n571), .B2(new_n291), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n569), .B(new_n570), .C1(new_n572), .C2(new_n358), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n573), .A2(KEYINPUT83), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(KEYINPUT83), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n309), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n574), .A2(new_n378), .A3(new_n575), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n291), .A2(new_n217), .A3(G68), .ZN(new_n579));
  INV_X1    g0379(.A(G87), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n580), .A2(new_n352), .A3(new_n465), .ZN(new_n581));
  OAI211_X1 g0381(.A(KEYINPUT19), .B(new_n581), .C1(new_n353), .C2(G20), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n254), .A2(new_n352), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n579), .B(new_n582), .C1(KEYINPUT19), .C2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n252), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n321), .A2(new_n328), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n464), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n327), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n577), .A2(new_n578), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n576), .A2(G190), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n574), .A2(G200), .A3(new_n575), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n585), .B(new_n586), .C1(new_n580), .C2(new_n464), .ZN(new_n595));
  INV_X1    g0395(.A(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n593), .A2(new_n594), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g0397(.A1(new_n592), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n565), .A2(KEYINPUT21), .A3(G169), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n309), .B2(new_n565), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n555), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n555), .A2(G169), .A3(new_n565), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT86), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT21), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n555), .A2(new_n565), .A3(KEYINPUT86), .A4(G169), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  AND2_X1   g0407(.A1(new_n486), .A2(G169), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n486), .A2(new_n309), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT88), .ZN(new_n610));
  OR3_X1    g0410(.A1(new_n608), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n610), .B1(new_n608), .B2(new_n609), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n598), .A2(new_n601), .A3(new_n607), .A4(new_n614), .ZN(new_n615));
  AND4_X1   g0415(.A1(new_n447), .A2(new_n544), .A3(new_n567), .A4(new_n615), .ZN(G372));
  NAND2_X1  g0416(.A1(new_n427), .A2(new_n428), .ZN(new_n617));
  AND3_X1   g0417(.A1(new_n443), .A2(KEYINPUT18), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(KEYINPUT18), .B1(new_n443), .B2(new_n617), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(new_n332), .ZN(new_n622));
  INV_X1    g0422(.A(new_n376), .ZN(new_n623));
  AOI22_X1  g0423(.A1(new_n383), .A2(new_n384), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n437), .A2(new_n440), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n621), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n626), .A2(new_n304), .A3(new_n308), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n627), .A2(new_n311), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n531), .A2(new_n536), .A3(new_n543), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n576), .A2(new_n309), .B1(new_n590), .B2(new_n588), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n573), .A2(new_n378), .ZN(new_n631));
  XOR2_X1   g0431(.A(new_n631), .B(KEYINPUT90), .Z(new_n632));
  AOI21_X1  g0432(.A(new_n595), .B1(new_n576), .B2(G190), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n573), .A2(G200), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n630), .A2(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OR2_X1    g0435(.A1(new_n608), .A2(new_n609), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n612), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n607), .A2(new_n601), .A3(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n629), .A2(new_n499), .A3(new_n635), .A4(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n536), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT26), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n640), .A2(new_n635), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n592), .A2(new_n597), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT26), .B1(new_n643), .B2(new_n536), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n630), .A2(new_n632), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n447), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n628), .A2(new_n648), .ZN(G369));
  NAND2_X1  g0449(.A1(new_n607), .A2(new_n601), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n229), .A2(G20), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n651), .A2(new_n216), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(G213), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g0455(.A(KEYINPUT91), .B(G343), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n556), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n650), .B(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n661), .A2(new_n567), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G330), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n499), .A2(new_n614), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n472), .B2(new_n659), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n614), .A2(new_n659), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n664), .A2(new_n650), .A3(new_n659), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n636), .A2(new_n612), .A3(new_n659), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g0474(.A(new_n674), .B(KEYINPUT92), .ZN(G399));
  INV_X1    g0475(.A(new_n231), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n676), .A2(G41), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n581), .A2(G116), .ZN(new_n678));
  NOR3_X1   g0478(.A1(new_n677), .A2(new_n216), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n679), .B1(new_n222), .B2(new_n677), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT28), .Z(new_n681));
  INV_X1    g0481(.A(KEYINPUT29), .ZN(new_n682));
  INV_X1    g0482(.A(new_n650), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n614), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n633), .A2(new_n634), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n544), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n598), .A2(new_n640), .A3(new_n641), .ZN(new_n687));
  AOI21_X1  g0487(.A(new_n641), .B1(new_n640), .B2(new_n635), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n688), .B1(new_n630), .B2(new_n632), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n686), .A2(new_n687), .A3(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n682), .B1(new_n690), .B2(new_n659), .ZN(new_n691));
  AOI211_X1 g0491(.A(KEYINPUT29), .B(new_n658), .C1(new_n639), .C2(new_n646), .ZN(new_n692));
  OR2_X1    g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n544), .A2(new_n615), .A3(new_n567), .A4(new_n659), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n524), .A2(new_n486), .A3(new_n309), .ZN(new_n695));
  INV_X1    g0495(.A(new_n564), .ZN(new_n696));
  AOI22_X1  g0496(.A1(new_n696), .A2(new_n562), .B1(G270), .B2(new_n484), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n695), .A2(new_n697), .A3(new_n576), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g0500(.A1(new_n573), .A2(new_n309), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n565), .A2(new_n701), .A3(new_n486), .A4(new_n524), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n695), .A2(KEYINPUT30), .A3(new_n697), .A4(new_n576), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n700), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT93), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n704), .A2(new_n658), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT31), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n706), .A3(new_n709), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n694), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n693), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n681), .B1(new_n716), .B2(G1), .ZN(G364));
  INV_X1    g0517(.A(new_n663), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n216), .B1(new_n651), .B2(G45), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n677), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n718), .A2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(G330), .B2(new_n662), .ZN(new_n723));
  INV_X1    g0523(.A(new_n721), .ZN(new_n724));
  XNOR2_X1  g0524(.A(KEYINPUT95), .B(G169), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n224), .B1(new_n725), .B2(G20), .ZN(new_n726));
  INV_X1    g0526(.A(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n334), .A2(new_n434), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n217), .A2(new_n309), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G326), .ZN(new_n732));
  INV_X1    g0532(.A(new_n729), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n733), .A2(new_n334), .A3(G200), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(G322), .ZN(new_n736));
  OAI211_X1 g0536(.A(new_n365), .B(new_n732), .C1(new_n735), .C2(new_n736), .ZN(new_n737));
  NOR3_X1   g0537(.A1(new_n733), .A2(new_n434), .A3(G190), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  XOR2_X1   g0539(.A(KEYINPUT33), .B(G317), .Z(new_n740));
  NOR3_X1   g0540(.A1(new_n733), .A2(G190), .A3(G200), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G311), .ZN(new_n743));
  OAI22_X1  g0543(.A1(new_n739), .A2(new_n740), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n728), .A2(G20), .A3(new_n309), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n737), .B(new_n744), .C1(G303), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n334), .A2(G20), .ZN(new_n748));
  XNOR2_X1  g0548(.A(new_n748), .B(KEYINPUT96), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n309), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n434), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(G200), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G283), .A2(new_n751), .B1(new_n752), .B2(G329), .ZN(new_n753));
  INV_X1    g0553(.A(G294), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n334), .A2(G179), .A3(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n217), .ZN(new_n756));
  OAI211_X1 g0556(.A(new_n747), .B(new_n753), .C1(new_n754), .C2(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n756), .A2(new_n352), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n746), .A2(G87), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n291), .B(new_n759), .C1(new_n735), .C2(new_n201), .ZN(new_n760));
  AOI211_X1 g0560(.A(new_n758), .B(new_n760), .C1(G50), .C2(new_n731), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n742), .A2(new_n322), .B1(new_n739), .B2(new_n202), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n751), .B2(G107), .ZN(new_n763));
  AOI21_X1  g0563(.A(KEYINPUT32), .B1(new_n752), .B2(G159), .ZN(new_n764));
  AND3_X1   g0564(.A1(new_n752), .A2(KEYINPUT32), .A3(G159), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n761), .B(new_n763), .C1(new_n764), .C2(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n727), .B1(new_n757), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT94), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n726), .ZN(new_n771));
  INV_X1    g0571(.A(new_n396), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n291), .A2(KEYINPUT75), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n676), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(new_n275), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n776), .B1(new_n223), .B2(new_n777), .C1(new_n287), .C2(new_n246), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n676), .A2(new_n365), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G355), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n778), .B(new_n780), .C1(G116), .C2(new_n231), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n767), .B1(new_n771), .B2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n770), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n782), .B1(new_n662), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n723), .B1(new_n724), .B2(new_n784), .ZN(G396));
  AOI21_X1  g0585(.A(new_n658), .B1(new_n639), .B2(new_n646), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n622), .A2(new_n658), .ZN(new_n787));
  INV_X1    g0587(.A(KEYINPUT100), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n787), .B(new_n788), .ZN(new_n789));
  AND2_X1   g0589(.A1(new_n331), .A2(new_n658), .ZN(new_n790));
  OR2_X1    g0590(.A1(new_n336), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g0592(.A(new_n786), .B(new_n792), .Z(new_n793));
  AOI21_X1  g0593(.A(new_n721), .B1(new_n793), .B2(new_n715), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n794), .A2(KEYINPUT101), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(KEYINPUT101), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n795), .B(new_n796), .C1(new_n715), .C2(new_n793), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n774), .B1(new_n752), .B2(G132), .ZN(new_n798));
  XOR2_X1   g0598(.A(new_n798), .B(KEYINPUT98), .Z(new_n799));
  INV_X1    g0599(.A(new_n751), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(new_n202), .ZN(new_n801));
  INV_X1    g0601(.A(new_n756), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n801), .B1(G58), .B2(new_n802), .ZN(new_n803));
  OAI211_X1 g0603(.A(new_n799), .B(new_n803), .C1(new_n212), .C2(new_n745), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n804), .B(KEYINPUT99), .Z(new_n805));
  AOI22_X1  g0605(.A1(G143), .A2(new_n734), .B1(new_n738), .B2(G150), .ZN(new_n806));
  INV_X1    g0606(.A(G137), .ZN(new_n807));
  INV_X1    g0607(.A(G159), .ZN(new_n808));
  OAI221_X1 g0608(.A(new_n806), .B1(new_n807), .B2(new_n730), .C1(new_n808), .C2(new_n742), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT34), .Z(new_n810));
  NOR2_X1   g0610(.A1(new_n805), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(G283), .ZN(new_n812));
  OR2_X1    g0612(.A1(new_n738), .A2(KEYINPUT97), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n738), .A2(KEYINPUT97), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI22_X1  g0615(.A1(new_n812), .A2(new_n815), .B1(new_n800), .B2(new_n580), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n745), .A2(new_n465), .ZN(new_n817));
  AOI211_X1 g0617(.A(new_n291), .B(new_n817), .C1(G294), .C2(new_n734), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n758), .B1(G116), .B2(new_n741), .ZN(new_n819));
  INV_X1    g0619(.A(new_n752), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n818), .B(new_n819), .C1(new_n820), .C2(new_n743), .ZN(new_n821));
  AOI211_X1 g0621(.A(new_n816), .B(new_n821), .C1(G303), .C2(new_n731), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n726), .B1(new_n811), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n823), .A2(new_n721), .ZN(new_n824));
  INV_X1    g0624(.A(new_n769), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n726), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n824), .B1(G77), .B2(new_n827), .C1(new_n769), .C2(new_n792), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n797), .A2(new_n828), .ZN(G384));
  NAND3_X1  g0629(.A1(new_n694), .A2(new_n710), .A3(new_n705), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n383), .A2(new_n384), .A3(new_n658), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT103), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n384), .A2(new_n658), .ZN(new_n833));
  AND3_X1   g0633(.A1(new_n385), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n832), .B1(new_n385), .B2(new_n833), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n830), .A2(new_n836), .A3(new_n792), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT38), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n442), .A2(new_n443), .ZN(new_n839));
  INV_X1    g0639(.A(new_n655), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n443), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT37), .ZN(new_n842));
  NAND4_X1  g0642(.A1(new_n839), .A2(new_n841), .A3(new_n842), .A4(new_n438), .ZN(new_n843));
  INV_X1    g0643(.A(new_n438), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT7), .B1(new_n774), .B2(new_n217), .ZN(new_n845));
  OAI21_X1  g0645(.A(G68), .B1(new_n845), .B2(new_n394), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT16), .B1(new_n846), .B2(new_n390), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n411), .B1(new_n847), .B2(new_n401), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n427), .A2(new_n428), .A3(new_n655), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(KEYINPUT37), .B1(new_n844), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n848), .A2(new_n840), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  AOI221_X4 g0653(.A(new_n838), .B1(new_n843), .B2(new_n851), .C1(new_n446), .C2(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n443), .B(new_n840), .C1(new_n620), .C2(new_n625), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n443), .A2(new_n849), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n856), .A2(KEYINPUT105), .A3(new_n438), .ZN(new_n857));
  OR2_X1    g0657(.A1(new_n438), .A2(KEYINPUT105), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n857), .A2(new_n858), .A3(KEYINPUT37), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(new_n843), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT38), .B1(new_n855), .B2(new_n860), .ZN(new_n861));
  OAI211_X1 g0661(.A(new_n837), .B(KEYINPUT40), .C1(new_n854), .C2(new_n861), .ZN(new_n862));
  AOI22_X1  g0662(.A1(new_n446), .A2(new_n853), .B1(new_n851), .B2(new_n843), .ZN(new_n863));
  OAI21_X1  g0663(.A(KEYINPUT104), .B1(new_n863), .B2(KEYINPUT38), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(KEYINPUT38), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT104), .ZN(new_n866));
  AND3_X1   g0666(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n444), .B1(new_n442), .B2(new_n443), .ZN(new_n868));
  NOR2_X1   g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  XNOR2_X1  g0669(.A(new_n438), .B(KEYINPUT17), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n852), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n843), .A2(new_n851), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n866), .B(new_n838), .C1(new_n871), .C2(new_n872), .ZN(new_n873));
  NAND3_X1  g0673(.A1(new_n864), .A2(new_n865), .A3(new_n873), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n874), .A2(new_n837), .ZN(new_n875));
  OAI211_X1 g0675(.A(G330), .B(new_n862), .C1(new_n875), .C2(KEYINPUT40), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n447), .A2(G330), .A3(new_n830), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g0678(.A(new_n878), .B(KEYINPUT107), .Z(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT40), .B1(new_n874), .B2(new_n837), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n861), .A2(new_n854), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n830), .A2(new_n836), .A3(new_n792), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT40), .ZN(new_n883));
  NOR3_X1   g0683(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n447), .A2(new_n830), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n879), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g0688(.A(new_n888), .B(KEYINPUT106), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n447), .B1(new_n691), .B2(new_n692), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n628), .ZN(new_n891));
  XNOR2_X1  g0691(.A(new_n889), .B(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n383), .A2(new_n384), .A3(new_n659), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT39), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n881), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n893), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n836), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n786), .A2(new_n792), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n332), .A2(new_n658), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n898), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g0702(.A1(new_n902), .A2(new_n874), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n621), .A2(new_n840), .ZN(new_n904));
  NOR3_X1   g0704(.A1(new_n897), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n892), .B(new_n905), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n216), .B2(new_n651), .ZN(new_n907));
  OAI211_X1 g0707(.A(G20), .B(new_n357), .C1(new_n506), .C2(KEYINPUT35), .ZN(new_n908));
  AOI211_X1 g0708(.A(new_n207), .B(new_n908), .C1(KEYINPUT35), .C2(new_n506), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT36), .Z(new_n910));
  OAI211_X1 g0710(.A(new_n222), .B(G77), .C1(new_n201), .C2(new_n202), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT102), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(G50), .B2(new_n202), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n913), .A2(G1), .A3(new_n229), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n907), .A2(new_n910), .A3(new_n914), .ZN(G367));
  NOR2_X1   g0715(.A1(new_n596), .A2(new_n659), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n635), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n645), .B2(new_n917), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n629), .B1(new_n541), .B2(new_n659), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n921), .A2(new_n671), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT42), .Z(new_n923));
  OR2_X1    g0723(.A1(new_n921), .A2(new_n614), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n658), .B1(new_n924), .B2(new_n536), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n920), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n919), .B(KEYINPUT108), .ZN(new_n927));
  XNOR2_X1  g0727(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n926), .B(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n921), .B1(new_n536), .B2(new_n659), .ZN(new_n931));
  AND2_X1   g0731(.A1(new_n669), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT110), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n930), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n932), .A2(new_n933), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n935), .B(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n716), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n673), .A2(new_n931), .ZN(new_n939));
  XNOR2_X1  g0739(.A(new_n939), .B(KEYINPUT44), .ZN(new_n940));
  INV_X1    g0740(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n673), .A2(new_n931), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT45), .ZN(new_n943));
  OAI211_X1 g0743(.A(KEYINPUT112), .B(new_n670), .C1(new_n941), .C2(new_n943), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n670), .A2(KEYINPUT112), .ZN(new_n945));
  INV_X1    g0745(.A(new_n943), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n670), .A2(KEYINPUT112), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .A4(new_n940), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n668), .B1(new_n683), .B2(new_n658), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT111), .ZN(new_n951));
  OR2_X1    g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n952), .A2(new_n671), .A3(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(new_n718), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n938), .B1(new_n949), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n677), .B(KEYINPUT41), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n719), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n937), .A2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n800), .A2(new_n322), .ZN(new_n961));
  INV_X1    g0761(.A(new_n815), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n961), .B1(G159), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n746), .A2(G58), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n752), .A2(G137), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n291), .B1(new_n735), .B2(new_n255), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n742), .A2(new_n212), .B1(new_n202), .B2(new_n756), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n966), .B(new_n967), .C1(G143), .C2(new_n731), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n963), .A2(new_n964), .A3(new_n965), .A4(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n774), .B1(new_n735), .B2(new_n558), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n746), .A2(KEYINPUT46), .A3(G116), .ZN(new_n971));
  OAI221_X1 g0771(.A(new_n971), .B1(new_n465), .B2(new_n756), .C1(new_n742), .C2(new_n812), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n970), .B(new_n972), .C1(G311), .C2(new_n731), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n962), .A2(G294), .B1(G97), .B2(new_n751), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n745), .A2(new_n207), .ZN(new_n975));
  OAI211_X1 g0775(.A(new_n973), .B(new_n974), .C1(KEYINPUT46), .C2(new_n975), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n752), .A2(G317), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n969), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT47), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n724), .B1(new_n979), .B2(new_n726), .ZN(new_n980));
  INV_X1    g0780(.A(new_n776), .ZN(new_n981));
  OAI221_X1 g0781(.A(new_n771), .B1(new_n231), .B2(new_n328), .C1(new_n981), .C2(new_n242), .ZN(new_n982));
  OAI211_X1 g0782(.A(new_n980), .B(new_n982), .C1(new_n783), .C2(new_n919), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n960), .A2(new_n983), .ZN(G387));
  AND2_X1   g0784(.A1(new_n752), .A2(G326), .ZN(new_n985));
  AOI22_X1  g0785(.A1(G303), .A2(new_n741), .B1(new_n734), .B2(G317), .ZN(new_n986));
  OAI221_X1 g0786(.A(new_n986), .B1(new_n736), .B2(new_n730), .C1(new_n815), .C2(new_n743), .ZN(new_n987));
  XNOR2_X1  g0787(.A(new_n987), .B(KEYINPUT48), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n812), .B2(new_n756), .C1(new_n754), .C2(new_n745), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT49), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n775), .B(new_n985), .C1(new_n989), .C2(new_n990), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n990), .B2(new_n989), .C1(new_n207), .C2(new_n800), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n735), .A2(new_n212), .B1(new_n322), .B2(new_n745), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n775), .B1(new_n742), .B2(new_n202), .C1(new_n253), .C2(new_n739), .ZN(new_n994));
  AOI211_X1 g0794(.A(new_n993), .B(new_n994), .C1(G159), .C2(new_n731), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n802), .A2(new_n327), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G97), .A2(new_n751), .B1(new_n752), .B2(G150), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n995), .A2(new_n996), .A3(new_n997), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n992), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n721), .B1(new_n999), .B2(new_n727), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n981), .B1(new_n239), .B2(new_n777), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n678), .B2(new_n779), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n253), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n1003), .B1(new_n1004), .B2(new_n212), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1005), .A2(new_n678), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1004), .A2(new_n1003), .A3(new_n212), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1006), .A2(new_n287), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g0808(.A(new_n1008), .B1(G68), .B2(G77), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n1002), .A2(new_n1009), .B1(G107), .B2(new_n231), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n1000), .B1(new_n771), .B2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n1011), .B(KEYINPUT114), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n667), .B2(new_n783), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n955), .A2(new_n720), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n955), .A2(new_n716), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n954), .B(new_n663), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n938), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1015), .A2(new_n1017), .A3(new_n677), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1013), .A2(new_n1014), .A3(new_n1018), .ZN(G393));
  OAI221_X1 g0819(.A(new_n771), .B1(new_n352), .B2(new_n231), .C1(new_n981), .C2(new_n249), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n775), .B1(new_n202), .B2(new_n745), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n734), .A2(G159), .B1(new_n731), .B2(G150), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT51), .ZN(new_n1023));
  AOI211_X1 g0823(.A(new_n1021), .B(new_n1023), .C1(new_n1004), .C2(new_n741), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n752), .A2(G143), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n802), .A2(G77), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n962), .A2(G50), .B1(G87), .B2(new_n751), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1024), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n365), .B1(new_n756), .B2(new_n207), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n734), .A2(G311), .B1(new_n731), .B2(G317), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT52), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(G294), .C2(new_n741), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(new_n962), .A2(G303), .B1(G107), .B2(new_n751), .ZN(new_n1033));
  OAI211_X1 g0833(.A(new_n1032), .B(new_n1033), .C1(new_n812), .C2(new_n745), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n820), .A2(new_n736), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1028), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n724), .B1(new_n1036), .B2(new_n726), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1020), .B(new_n1037), .C1(new_n931), .C2(new_n783), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n949), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1038), .B1(new_n1039), .B2(new_n719), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n677), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n1039), .B2(new_n1015), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n955), .A2(new_n949), .A3(new_n716), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1040), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(G390));
  AOI21_X1  g0845(.A(new_n900), .B1(new_n786), .B2(new_n792), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n893), .B1(new_n1046), .B2(new_n898), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n894), .A2(new_n1047), .A3(new_n896), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n690), .A2(new_n659), .A3(new_n792), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n901), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1050), .A2(new_n836), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n893), .B(KEYINPUT115), .Z(new_n1052));
  NOR2_X1   g0852(.A1(new_n881), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(G330), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n789), .B2(new_n791), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n713), .A2(new_n836), .A3(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n1048), .A2(new_n1054), .A3(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(KEYINPUT117), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1048), .A2(new_n1054), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n830), .A2(new_n836), .A3(new_n1056), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(KEYINPUT116), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT116), .ZN(new_n1063));
  NAND4_X1  g0863(.A1(new_n830), .A2(new_n836), .A3(new_n1063), .A4(new_n1056), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1060), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(KEYINPUT117), .ZN(new_n1067));
  NAND4_X1  g0867(.A1(new_n1048), .A2(new_n1054), .A3(new_n1067), .A4(new_n1057), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1059), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  OR2_X1    g0869(.A1(new_n1069), .A2(new_n719), .ZN(new_n1070));
  NOR3_X1   g0870(.A1(new_n861), .A2(new_n854), .A3(KEYINPUT39), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(KEYINPUT39), .B2(new_n874), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n825), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n962), .A2(G107), .B1(G97), .B2(new_n741), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n1074), .B1(new_n812), .B2(new_n730), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT119), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n365), .B(new_n1026), .C1(new_n735), .C2(new_n207), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(new_n752), .B2(G294), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1077), .A2(new_n759), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1081));
  NOR3_X1   g0881(.A1(new_n745), .A2(KEYINPUT53), .A3(new_n255), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n291), .B1(new_n800), .B2(new_n212), .ZN(new_n1083));
  OR2_X1    g0883(.A1(new_n1083), .A2(KEYINPUT118), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(KEYINPUT118), .ZN(new_n1085));
  AOI22_X1  g0885(.A1(new_n962), .A2(G137), .B1(G125), .B2(new_n752), .ZN(new_n1086));
  OAI21_X1  g0886(.A(KEYINPUT53), .B1(new_n745), .B2(new_n255), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n808), .B2(new_n756), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n734), .A2(G132), .ZN(new_n1089));
  XOR2_X1   g0889(.A(KEYINPUT54), .B(G143), .Z(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1089), .B1(new_n742), .B2(new_n1091), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1088), .B(new_n1092), .C1(G128), .C2(new_n731), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1084), .A2(new_n1085), .A3(new_n1086), .A4(new_n1093), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1081), .A2(new_n801), .B1(new_n1082), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n724), .B1(new_n1095), .B2(new_n726), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1073), .B(new_n1096), .C1(new_n1004), .C2(new_n827), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n890), .A2(new_n628), .A3(new_n877), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n713), .A2(new_n1056), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n898), .ZN(new_n1100));
  NAND3_X1  g0900(.A1(new_n1062), .A2(new_n1064), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1046), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n830), .A2(new_n1056), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n898), .ZN(new_n1105));
  NAND4_X1  g0905(.A1(new_n1105), .A2(new_n901), .A3(new_n1049), .A4(new_n1057), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1098), .B1(new_n1103), .B2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  AND2_X1   g0908(.A1(new_n1069), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1059), .A2(new_n1066), .A3(new_n1068), .A4(new_n1107), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(new_n677), .ZN(new_n1111));
  OAI211_X1 g0911(.A(new_n1070), .B(new_n1097), .C1(new_n1109), .C2(new_n1111), .ZN(G378));
  INV_X1    g0912(.A(new_n904), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n902), .A2(new_n874), .ZN(new_n1114));
  OAI211_X1 g0914(.A(new_n1113), .B(new_n1114), .C1(new_n1072), .C2(new_n893), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(KEYINPUT120), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n312), .A2(KEYINPUT55), .ZN(new_n1117));
  INV_X1    g0917(.A(KEYINPUT55), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n304), .A2(new_n308), .A3(new_n1118), .A4(new_n311), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n269), .A2(new_n840), .ZN(new_n1120));
  XOR2_X1   g0920(.A(new_n1120), .B(KEYINPUT56), .Z(new_n1121));
  AND3_X1   g0921(.A1(new_n1117), .A2(new_n1119), .A3(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1121), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n885), .B2(G330), .ZN(new_n1126));
  NOR4_X1   g0926(.A1(new_n880), .A2(new_n884), .A3(new_n1055), .A4(new_n1124), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1116), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n876), .A2(new_n1124), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n885), .A2(G330), .A3(new_n1125), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1129), .A2(new_n1130), .A3(KEYINPUT120), .A4(new_n1115), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1128), .A2(new_n720), .A3(new_n1131), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n276), .B1(new_n322), .B2(new_n745), .C1(new_n735), .C2(new_n465), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n774), .B1(new_n202), .B2(new_n756), .C1(new_n742), .C2(new_n328), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(G116), .C2(new_n731), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(G58), .A2(new_n751), .B1(new_n752), .B2(G283), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1135), .B(new_n1136), .C1(new_n352), .C2(new_n739), .ZN(new_n1137));
  XNOR2_X1  g0937(.A(new_n1137), .B(KEYINPUT58), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n742), .A2(new_n807), .B1(new_n255), .B2(new_n756), .ZN(new_n1139));
  AOI22_X1  g0939(.A1(new_n734), .A2(G128), .B1(new_n731), .B2(G125), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n745), .B2(new_n1091), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1139), .B(new_n1141), .C1(G132), .C2(new_n738), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT59), .ZN(new_n1143));
  AOI21_X1  g0943(.A(G41), .B1(new_n752), .B2(G124), .ZN(new_n1144));
  AOI21_X1  g0944(.A(G33), .B1(new_n751), .B2(G159), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n1144), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(G41), .B1(new_n775), .B2(G33), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1138), .B(new_n1146), .C1(G50), .C2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n724), .B1(new_n1148), .B2(new_n726), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1149), .B1(G50), .B2(new_n827), .C1(new_n1125), .C2(new_n769), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1132), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT57), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1098), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1110), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1152), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1115), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1129), .A2(new_n905), .A3(new_n1130), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n1152), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1110), .A2(new_n1153), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1041), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1151), .B1(new_n1156), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(G375));
  NOR2_X1   g0963(.A1(new_n836), .A2(new_n769), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n827), .A2(G68), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n291), .B1(new_n731), .B2(G294), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1166), .B(new_n996), .C1(new_n742), .C2(new_n465), .ZN(new_n1167));
  NOR2_X1   g0967(.A1(new_n961), .A2(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1168), .B1(new_n207), .B2(new_n815), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n820), .A2(new_n558), .B1(new_n352), .B2(new_n745), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1169), .B1(KEYINPUT122), .B2(new_n1170), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(KEYINPUT122), .B2(new_n1170), .C1(new_n812), .C2(new_n735), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(G159), .A2(new_n746), .B1(new_n731), .B2(G132), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1173), .B1(new_n807), .B2(new_n735), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n774), .B(new_n1174), .C1(G150), .C2(new_n741), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n752), .A2(G128), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n802), .A2(G50), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n962), .A2(new_n1090), .B1(G58), .B2(new_n751), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .A4(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n727), .B1(new_n1172), .B2(new_n1179), .ZN(new_n1180));
  NOR4_X1   g0980(.A1(new_n1164), .A2(new_n724), .A3(new_n1165), .A4(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n719), .B(KEYINPUT121), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1181), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1103), .A2(new_n1098), .A3(new_n1106), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n957), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1184), .B1(new_n1186), .B2(new_n1107), .ZN(G381));
  INV_X1    g0987(.A(G378), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1162), .A2(new_n1188), .ZN(new_n1189));
  NOR3_X1   g0989(.A1(new_n1189), .A2(G384), .A3(G381), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n960), .A2(new_n1044), .A3(new_n983), .ZN(new_n1191));
  INV_X1    g0991(.A(new_n1191), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(G393), .A2(G396), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n1190), .A2(new_n1192), .A3(new_n1193), .ZN(G407));
  OAI211_X1 g0994(.A(G407), .B(G213), .C1(new_n656), .C2(new_n1189), .ZN(G409));
  NAND2_X1  g0995(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n1183), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n1150), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(KEYINPUT124), .ZN(new_n1199));
  NOR3_X1   g0999(.A1(new_n1116), .A2(new_n1126), .A3(new_n1127), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n1129), .A2(new_n1130), .B1(new_n1115), .B2(KEYINPUT120), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1202), .A2(new_n957), .A3(new_n1160), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT124), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1197), .A2(new_n1204), .A3(new_n1150), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1199), .A2(new_n1203), .A3(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1206), .A2(new_n1188), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1151), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(new_n677), .ZN(new_n1210));
  AOI21_X1  g1010(.A(KEYINPUT57), .B1(new_n1202), .B2(new_n1160), .ZN(new_n1211));
  OAI211_X1 g1011(.A(G378), .B(new_n1208), .C1(new_n1210), .C2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT123), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  AOI21_X1  g1014(.A(KEYINPUT123), .B1(new_n1162), .B2(G378), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1207), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n657), .A2(G213), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT60), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1107), .B1(new_n1218), .B2(new_n1185), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n677), .C1(new_n1218), .C2(new_n1185), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1220), .A2(new_n1184), .ZN(new_n1221));
  AND2_X1   g1021(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1221), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1216), .A2(new_n1217), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(KEYINPUT62), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT61), .ZN(new_n1230));
  INV_X1    g1030(.A(G2897), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1226), .B1(new_n1231), .B2(new_n1217), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1217), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1223), .A2(G2897), .A3(new_n1233), .A4(new_n1225), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1232), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1162), .A2(KEYINPUT123), .A3(G378), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n1236), .A2(new_n1237), .B1(new_n1188), .B2(new_n1206), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1235), .B1(new_n1238), .B2(new_n1233), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT62), .ZN(new_n1240));
  NAND4_X1  g1040(.A1(new_n1216), .A2(new_n1240), .A3(new_n1217), .A4(new_n1227), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1229), .A2(new_n1230), .A3(new_n1239), .A4(new_n1241), .ZN(new_n1242));
  AND2_X1   g1042(.A1(G393), .A2(G396), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1243), .A2(new_n1193), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1044), .B1(new_n960), .B2(new_n983), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1244), .B1(new_n1192), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1245), .ZN(new_n1247));
  XNOR2_X1  g1047(.A(G393), .B(G396), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(new_n1248), .A3(new_n1191), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1246), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1242), .A2(new_n1250), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n1238), .A2(new_n1233), .A3(new_n1226), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT126), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1246), .A2(new_n1249), .A3(new_n1230), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n1252), .A2(KEYINPUT63), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  AOI22_X1  g1055(.A1(new_n1216), .A2(new_n1217), .B1(new_n1232), .B2(new_n1234), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT63), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1228), .B1(new_n1256), .B2(new_n1257), .ZN(new_n1258));
  OR2_X1    g1058(.A1(new_n1254), .A2(new_n1253), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1255), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1251), .A2(new_n1260), .ZN(G405));
  OR2_X1    g1061(.A1(new_n1226), .A2(KEYINPUT127), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1250), .B(new_n1262), .ZN(new_n1263));
  AOI22_X1  g1063(.A1(new_n1236), .A2(new_n1237), .B1(new_n1188), .B2(G375), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1263), .B(new_n1264), .ZN(G402));
endmodule


